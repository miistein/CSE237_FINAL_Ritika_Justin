module conv7 (
input clock,
input reset,
input vld_in,
input [191:0][0:0] in,
output vld_out,
output [63:0][0:0] out
);
reg [6:0] vld_reg = 0;
wire [6:0] resets;
reg [5:0] rst_reg;
assign resets = { rst_reg, reset };
assign vld_out = vld_reg[6];
always @( posedge clock ) begin
vld_reg <= { vld_reg[5:0], vld_in };
rst_reg <= resets[5:0];
end
wire [0:0] tree_0;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_192 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[111]),
 .b(in[158]),
 .c(tree_0)
);
wire [0:0] tree_1;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_193 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[56]),
 .b(in[130]),
 .c(tree_1)
);
wire [0:0] tree_2;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_194 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[118]),
 .b(in[161]),
 .c(tree_2)
);
wire [0:0] tree_3;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_195 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[125]),
 .b(in[182]),
 .c(tree_3)
);
wire [0:0] tree_4;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_196 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[38]),
 .b(in[179]),
 .c(tree_4)
);
wire [0:0] tree_5;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_197 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[74]),
 .b(in[83]),
 .c(tree_5)
);
wire [0:0] tree_6;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_198 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[36]),
 .b(in[175]),
 .c(tree_6)
);
wire [0:0] tree_7;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_199 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[46]),
 .b(in[99]),
 .c(tree_7)
);
wire [0:0] tree_8;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_200 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[80]),
 .b(in[178]),
 .c(tree_8)
);
wire [0:0] tree_9;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_201 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[17]),
 .b(in[66]),
 .c(tree_9)
);
wire [0:0] tree_10;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_202 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[19]),
 .b(in[133]),
 .c(tree_10)
);
wire [0:0] tree_11;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_203 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[82]),
 .b(in[155]),
 .c(tree_11)
);
wire [0:0] tree_12;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_204 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[97]),
 .b(in[140]),
 .c(tree_12)
);
wire [0:0] tree_13;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_205 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[124]),
 .b(in[183]),
 .c(tree_13)
);
wire [0:0] tree_14;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_206 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[63]),
 .b(in[166]),
 .c(tree_14)
);
wire [0:0] tree_15;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_207 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[12]),
 .b(in[44]),
 .c(tree_15)
);
wire [0:0] tree_16;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_208 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[55]),
 .b(in[170]),
 .c(tree_16)
);
wire [0:0] tree_17;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_209 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[39]),
 .b(in[105]),
 .c(tree_17)
);
wire [0:0] tree_18;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_210 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[95]),
 .b(in[167]),
 .c(tree_18)
);
wire [0:0] tree_19;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_211 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[20]),
 .b(in[48]),
 .c(tree_19)
);
wire [0:0] tree_20;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_212 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[148]),
 .b(in[188]),
 .c(tree_20)
);
wire [0:0] tree_21;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_213 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[21]),
 .b(in[47]),
 .c(tree_21)
);
wire [0:0] tree_22;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_214 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[53]),
 .b(in[119]),
 .c(tree_22)
);
wire [0:0] tree_23;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_215 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[27]),
 .b(in[173]),
 .c(tree_23)
);
wire [0:0] tree_24;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_216 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[151]),
 .b(in[168]),
 .c(tree_24)
);
wire [0:0] tree_25;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_217 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[77]),
 .b(in[181]),
 .c(tree_25)
);
wire [0:0] tree_26;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_218 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[24]),
 .b(in[163]),
 .c(tree_26)
);
wire [0:0] tree_27;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_219 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[7]),
 .b(in[9]),
 .c(tree_27)
);
wire [0:0] tree_28;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_220 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[87]),
 .b(in[156]),
 .c(tree_28)
);
wire [0:0] tree_29;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_221 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[150]),
 .b(in[162]),
 .c(tree_29)
);
wire [0:0] tree_30;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_222 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[5]),
 .b(in[94]),
 .c(tree_30)
);
wire [0:0] tree_31;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_223 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[71]),
 .b(in[131]),
 .c(tree_31)
);
wire [0:0] tree_32;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_224 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[11]),
 .b(in[162]),
 .c(tree_32)
);
wire [0:0] tree_33;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_225 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[80]),
 .b(in[135]),
 .c(tree_33)
);
wire [0:0] tree_34;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_226 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[3]),
 .b(in[79]),
 .c(tree_34)
);
wire [0:0] tree_35;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_227 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[54]),
 .b(in[112]),
 .c(tree_35)
);
wire [0:0] tree_36;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_228 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[77]),
 .b(in[182]),
 .c(tree_36)
);
wire [0:0] tree_37;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_229 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[86]),
 .b(in[122]),
 .c(tree_37)
);
wire [0:0] tree_38;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_230 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[27]),
 .b(in[134]),
 .c(tree_38)
);
wire [0:0] tree_39;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_231 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[2]),
 .b(in[178]),
 .c(tree_39)
);
wire [0:0] tree_40;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_232 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[124]),
 .b(in[169]),
 .c(tree_40)
);
wire [0:0] tree_41;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_233 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[40]),
 .b(in[109]),
 .c(tree_41)
);
wire [0:0] tree_42;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_234 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[36]),
 .b(in[71]),
 .c(tree_42)
);
wire [0:0] tree_43;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_235 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[81]),
 .b(in[95]),
 .c(tree_43)
);
wire [0:0] tree_44;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_236 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[102]),
 .b(in[188]),
 .c(tree_44)
);
wire [0:0] tree_45;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_237 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[89]),
 .b(in[107]),
 .c(tree_45)
);
wire [0:0] tree_46;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_238 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[39]),
 .b(in[103]),
 .c(tree_46)
);
wire [0:0] tree_47;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_239 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[5]),
 .b(in[37]),
 .c(tree_47)
);
wire [0:0] tree_48;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_240 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[7]),
 .b(in[16]),
 .c(tree_48)
);
wire [0:0] tree_49;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_241 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[66]),
 .b(in[116]),
 .c(tree_49)
);
wire [0:0] tree_50;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_242 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[0]),
 .b(in[100]),
 .c(tree_50)
);
wire [0:0] tree_51;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_243 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[31]),
 .b(in[57]),
 .c(tree_51)
);
wire [0:0] tree_52;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_244 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[65]),
 .b(in[160]),
 .c(tree_52)
);
wire [0:0] tree_53;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_245 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[59]),
 .b(in[91]),
 .c(tree_53)
);
wire [0:0] tree_54;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_246 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[22]),
 .b(in[145]),
 .c(tree_54)
);
wire [0:0] tree_55;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_247 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[4]),
 .b(in[30]),
 .c(tree_55)
);
wire [0:0] tree_56;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_248 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[24]),
 .b(in[104]),
 .c(tree_56)
);
wire [0:0] tree_57;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_249 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[90]),
 .b(in[115]),
 .c(tree_57)
);
wire [0:0] tree_58;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_250 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[43]),
 .b(in[60]),
 .c(tree_58)
);
wire [0:0] tree_59;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_251 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[41]),
 .b(in[131]),
 .c(tree_59)
);
wire [0:0] tree_60;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_252 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[28]),
 .b(in[48]),
 .c(tree_60)
);
wire [0:0] tree_61;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_253 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[52]),
 .b(in[180]),
 .c(tree_61)
);
wire [0:0] tree_62;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_254 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[37]),
 .b(in[174]),
 .c(tree_62)
);
wire [0:0] tree_63;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_255 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[92]),
 .b(in[112]),
 .c(tree_63)
);
wire [0:0] tree_64;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_256 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[19]),
 .b(in[120]),
 .c(tree_64)
);
wire [0:0] tree_65;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_257 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[39]),
 .b(in[116]),
 .c(tree_65)
);
wire [0:0] tree_66;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_258 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[59]),
 .b(in[167]),
 .c(tree_66)
);
wire [0:0] tree_67;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_259 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[101]),
 .b(in[190]),
 .c(tree_67)
);
wire [0:0] tree_68;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_260 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[146]),
 .b(in[153]),
 .c(tree_68)
);
wire [0:0] tree_69;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_261 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[16]),
 .b(in[18]),
 .c(tree_69)
);
wire [0:0] tree_70;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_262 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[70]),
 .b(in[137]),
 .c(tree_70)
);
wire [0:0] tree_71;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_263 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[30]),
 .b(in[128]),
 .c(tree_71)
);
wire [0:0] tree_72;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_264 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[33]),
 .b(in[94]),
 .c(tree_72)
);
wire [0:0] tree_73;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_265 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[157]),
 .b(in[176]),
 .c(tree_73)
);
wire [0:0] tree_74;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_266 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[12]),
 .b(in[90]),
 .c(tree_74)
);
wire [0:0] tree_75;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_267 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[126]),
 .b(in[130]),
 .c(tree_75)
);
wire [0:0] tree_76;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_268 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[144]),
 .b(in[185]),
 .c(tree_76)
);
wire [0:0] tree_77;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_269 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[6]),
 .b(in[149]),
 .c(tree_77)
);
wire [0:0] tree_78;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_270 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[50]),
 .b(in[187]),
 .c(tree_78)
);
wire [0:0] tree_79;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_271 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[51]),
 .b(in[115]),
 .c(tree_79)
);
wire [0:0] tree_80;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_272 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[94]),
 .b(in[191]),
 .c(tree_80)
);
wire [0:0] tree_81;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_273 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[91]),
 .b(in[173]),
 .c(tree_81)
);
wire [0:0] tree_82;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_274 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[77]),
 .b(in[104]),
 .c(tree_82)
);
wire [0:0] tree_83;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_275 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[70]),
 .b(in[105]),
 .c(tree_83)
);
wire [0:0] tree_84;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_276 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[49]),
 .b(in[169]),
 .c(tree_84)
);
wire [0:0] tree_85;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_277 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[146]),
 .b(in[147]),
 .c(tree_85)
);
wire [0:0] tree_86;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_278 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[35]),
 .b(in[189]),
 .c(tree_86)
);
wire [0:0] tree_87;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_279 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[62]),
 .b(in[93]),
 .c(tree_87)
);
wire [0:0] tree_88;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_280 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[101]),
 .b(in[171]),
 .c(tree_88)
);
wire [0:0] tree_89;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_281 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[21]),
 .b(in[142]),
 .c(tree_89)
);
wire [0:0] tree_90;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_282 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[108]),
 .b(in[170]),
 .c(tree_90)
);
wire [0:0] tree_91;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_283 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[85]),
 .b(in[153]),
 .c(tree_91)
);
wire [0:0] tree_92;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_284 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[135]),
 .b(1'h0),
 .c(tree_92)
);
wire [0:0] tree_93;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_285 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_92),
 .b(tree_37),
 .c(tree_93)
);
wire [0:0] tree_94;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_286 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[163]),
 .b(1'h0),
 .c(tree_94)
);
wire [0:0] tree_95;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_287 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_94),
 .b(tree_78),
 .c(tree_95)
);
wire [0:0] tree_96;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_288 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[8]),
 .b(in[80]),
 .c(tree_96)
);
wire [0:0] tree_97;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_289 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[34]),
 .b(in[69]),
 .c(tree_97)
);
wire [0:0] tree_98;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_290 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[20]),
 .b(in[112]),
 .c(tree_98)
);
wire [0:0] tree_99;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_291 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[48]),
 .b(in[127]),
 .c(tree_99)
);
wire [0:0] tree_100;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_292 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[19]),
 .b(in[88]),
 .c(tree_100)
);
wire [0:0] tree_101;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_293 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[32]),
 .b(in[126]),
 .c(tree_101)
);
wire [0:0] tree_102;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_294 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[46]),
 .b(in[52]),
 .c(tree_102)
);
wire [0:0] tree_103;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_295 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[84]),
 .b(in[129]),
 .c(tree_103)
);
wire [0:0] tree_104;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_296 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[86]),
 .b(in[184]),
 .c(tree_104)
);
wire [0:0] tree_105;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_297 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[22]),
 .b(in[159]),
 .c(tree_105)
);
wire [0:0] tree_106;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_298 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[121]),
 .b(in[122]),
 .c(tree_106)
);
wire [0:0] tree_107;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_299 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[67]),
 .b(in[90]),
 .c(tree_107)
);
wire [0:0] tree_108;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_300 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[26]),
 .b(in[89]),
 .c(tree_108)
);
wire [0:0] tree_109;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_301 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[102]),
 .b(1'h0),
 .c(tree_109)
);
wire [0:0] tree_110;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_302 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_109),
 .b(tree_84),
 .c(tree_110)
);
wire [0:0] tree_111;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_303 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[104]),
 .b(in[142]),
 .c(tree_111)
);
wire [0:0] tree_112;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_304 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[83]),
 .b(in[148]),
 .c(tree_112)
);
wire [0:0] tree_113;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_305 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[93]),
 .b(in[136]),
 .c(tree_113)
);
wire [0:0] tree_114;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_306 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[110]),
 .b(in[134]),
 .c(tree_114)
);
wire [0:0] tree_115;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_307 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[64]),
 .b(1'h0),
 .c(tree_115)
);
wire [0:0] tree_116;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_308 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_115),
 .b(tree_79),
 .c(tree_116)
);
wire [0:0] tree_117;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_309 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[133]),
 .b(in[181]),
 .c(tree_117)
);
wire [0:0] tree_118;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_310 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[25]),
 .b(in[149]),
 .c(tree_118)
);
wire [0:0] tree_119;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_311 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[103]),
 .b(in[175]),
 .c(tree_119)
);
wire [0:0] tree_120;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_312 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[45]),
 .b(in[160]),
 .c(tree_120)
);
wire [0:0] tree_121;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_313 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[11]),
 .b(in[41]),
 .c(tree_121)
);
wire [0:0] tree_122;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_314 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[78]),
 .b(in[86]),
 .c(tree_122)
);
wire [0:0] tree_123;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_315 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[98]),
 .b(in[119]),
 .c(tree_123)
);
wire [0:0] tree_124;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_316 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[29]),
 .b(in[122]),
 .c(tree_124)
);
wire [0:0] tree_125;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_317 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[39]),
 .b(in[49]),
 .c(tree_125)
);
wire [0:0] tree_126;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_318 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[84]),
 .b(in[106]),
 .c(tree_126)
);
wire [0:0] tree_127;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_319 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[128]),
 .b(1'h0),
 .c(tree_127)
);
wire [0:0] tree_128;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_320 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_127),
 .b(tree_26),
 .c(tree_128)
);
wire [0:0] tree_129;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_321 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[32]),
 .b(in[166]),
 .c(tree_129)
);
wire [0:0] tree_130;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_322 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[153]),
 .b(1'h0),
 .c(tree_130)
);
wire [0:0] tree_131;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_323 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_130),
 .b(tree_85),
 .c(tree_131)
);
wire [0:0] tree_132;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_324 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[62]),
 .b(in[97]),
 .c(tree_132)
);
wire [0:0] tree_133;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_325 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[88]),
 .b(in[168]),
 .c(tree_133)
);
wire [0:0] tree_134;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_326 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[89]),
 .b(in[154]),
 .c(tree_134)
);
wire [0:0] tree_135;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_327 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[90]),
 .b(in[141]),
 .c(tree_135)
);
wire [0:0] tree_136;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_328 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[35]),
 .b(in[138]),
 .c(tree_136)
);
wire [0:0] tree_137;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_329 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[43]),
 .b(in[60]),
 .c(tree_137)
);
wire [0:0] tree_138;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_330 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[73]),
 .b(in[76]),
 .c(tree_138)
);
wire [0:0] tree_139;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_331 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[113]),
 .b(in[177]),
 .c(tree_139)
);
wire [0:0] tree_140;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_332 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[8]),
 .b(in[190]),
 .c(tree_140)
);
wire [0:0] tree_141;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_333 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[48]),
 .b(in[125]),
 .c(tree_141)
);
wire [0:0] tree_142;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_334 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[180]),
 .b(1'h0),
 .c(tree_142)
);
wire [0:0] tree_143;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_335 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_142),
 .b(tree_6),
 .c(tree_143)
);
wire [0:0] tree_144;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_336 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[4]),
 .b(in[34]),
 .c(tree_144)
);
wire [0:0] tree_145;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_337 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[42]),
 .b(in[66]),
 .c(tree_145)
);
wire [0:0] tree_146;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_338 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[118]),
 .b(in[164]),
 .c(tree_146)
);
wire [0:0] tree_147;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_339 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[15]),
 .b(in[83]),
 .c(tree_147)
);
wire [0:0] tree_148;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_340 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[101]),
 .b(1'h0),
 .c(tree_148)
);
wire [0:0] tree_149;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_341 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_148),
 .b(tree_50),
 .c(tree_149)
);
wire [0:0] tree_150;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_342 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[135]),
 .b(in[143]),
 .c(tree_150)
);
wire [0:0] tree_151;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_343 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[97]),
 .b(in[159]),
 .c(tree_151)
);
wire [0:0] tree_152;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_344 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[147]),
 .b(in[182]),
 .c(tree_152)
);
wire [0:0] tree_153;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_345 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[82]),
 .b(in[105]),
 .c(tree_153)
);
wire [0:0] tree_154;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_346 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_30),
 .b(tree_107),
 .c(tree_154)
);
wire [0:0] tree_155;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_347 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[40]),
 .b(in[141]),
 .c(tree_155)
);
wire [0:0] tree_156;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_348 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[15]),
 .b(in[160]),
 .c(tree_156)
);
wire [0:0] tree_157;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_349 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[18]),
 .b(in[172]),
 .c(tree_157)
);
wire [0:0] tree_158;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_350 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[58]),
 .b(in[180]),
 .c(tree_158)
);
wire [0:0] tree_159;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_351 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[23]),
 .b(in[171]),
 .c(tree_159)
);
wire [0:0] tree_160;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_352 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[61]),
 .b(in[151]),
 .c(tree_160)
);
wire [0:0] tree_161;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_353 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[19]),
 .b(in[72]),
 .c(tree_161)
);
wire [0:0] tree_162;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_354 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[17]),
 .b(in[22]),
 .c(tree_162)
);
wire [0:0] tree_163;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_355 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[62]),
 .b(in[92]),
 .c(tree_163)
);
wire [0:0] tree_164;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_356 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[36]),
 .b(in[165]),
 .c(tree_164)
);
wire [0:0] tree_165;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_357 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[106]),
 .b(in[183]),
 .c(tree_165)
);
wire [0:0] tree_166;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_358 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[107]),
 .b(in[117]),
 .c(tree_166)
);
wire [0:0] tree_167;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_359 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[52]),
 .b(in[76]),
 .c(tree_167)
);
wire [0:0] tree_168;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_360 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[137]),
 .b(in[138]),
 .c(tree_168)
);
wire [0:0] tree_169;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_361 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[6]),
 .b(in[30]),
 .c(tree_169)
);
wire [0:0] tree_170;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_362 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[99]),
 .b(in[134]),
 .c(tree_170)
);
wire [0:0] tree_171;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_363 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[4]),
 .b(in[140]),
 .c(tree_171)
);
wire [0:0] tree_172;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_364 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[150]),
 .b(in[188]),
 .c(tree_172)
);
wire [0:0] tree_173;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_365 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[108]),
 .b(in[152]),
 .c(tree_173)
);
wire [0:0] tree_174;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_366 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[168]),
 .b(1'h0),
 .c(tree_174)
);
wire [0:0] tree_175;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_367 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_174),
 .b(tree_15),
 .c(tree_175)
);
wire [0:0] tree_176;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_368 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_49),
 .b(tree_166),
 .c(tree_176)
);
wire [0:0] tree_177;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_369 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_99),
 .b(tree_79),
 .c(tree_177)
);
wire [0:0] tree_178;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_370 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[97]),
 .b(1'h0),
 .c(tree_178)
);
wire [0:0] tree_179;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_371 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_178),
 .b(tree_27),
 .c(tree_179)
);
wire [0:0] tree_180;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_372 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[29]),
 .b(in[47]),
 .c(tree_180)
);
wire [0:0] tree_181;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_373 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[109]),
 .b(in[183]),
 .c(tree_181)
);
wire [0:0] tree_182;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_374 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[24]),
 .b(in[67]),
 .c(tree_182)
);
wire [0:0] tree_183;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_375 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[68]),
 .b(in[175]),
 .c(tree_183)
);
wire [0:0] tree_184;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_376 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[64]),
 .b(in[170]),
 .c(tree_184)
);
wire [0:0] tree_185;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_377 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[114]),
 .b(in[120]),
 .c(tree_185)
);
wire [0:0] tree_186;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_378 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[129]),
 .b(1'h0),
 .c(tree_186)
);
wire [0:0] tree_187;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_379 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_186),
 .b(tree_1),
 .c(tree_187)
);
wire [0:0] tree_188;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_380 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[102]),
 .b(in[135]),
 .c(tree_188)
);
wire [0:0] tree_189;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_381 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[3]),
 .b(in[33]),
 .c(tree_189)
);
wire [0:0] tree_190;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_382 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[39]),
 .b(in[132]),
 .c(tree_190)
);
wire [0:0] tree_191;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_383 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[2]),
 .b(in[171]),
 .c(tree_191)
);
wire [0:0] tree_192;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_384 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[54]),
 .b(in[80]),
 .c(tree_192)
);
wire [0:0] tree_193;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_385 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[5]),
 .b(in[164]),
 .c(tree_193)
);
wire [0:0] tree_194;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_386 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[37]),
 .b(in[123]),
 .c(tree_194)
);
wire [0:0] tree_195;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_387 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[91]),
 .b(in[96]),
 .c(tree_195)
);
wire [0:0] tree_196;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_388 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[98]),
 .b(1'h0),
 .c(tree_196)
);
wire [0:0] tree_197;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_389 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_196),
 .b(tree_181),
 .c(tree_197)
);
wire [0:0] tree_198;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_390 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[0]),
 .b(in[60]),
 .c(tree_198)
);
wire [0:0] tree_199;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_391 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[186]),
 .b(1'h0),
 .c(tree_199)
);
wire [0:0] tree_200;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_392 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_199),
 .b(tree_76),
 .c(tree_200)
);
wire [0:0] tree_201;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_393 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[51]),
 .b(in[85]),
 .c(tree_201)
);
wire [0:0] tree_202;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_394 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[107]),
 .b(in[148]),
 .c(tree_202)
);
wire [0:0] tree_203;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_395 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[28]),
 .b(1'h0),
 .c(tree_203)
);
wire [0:0] tree_204;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_396 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_203),
 .b(tree_139),
 .c(tree_204)
);
wire [0:0] tree_205;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_397 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[14]),
 .b(in[64]),
 .c(tree_205)
);
wire [0:0] tree_206;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_398 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[75]),
 .b(in[95]),
 .c(tree_206)
);
wire [0:0] tree_207;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_399 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[93]),
 .b(1'h0),
 .c(tree_207)
);
wire [0:0] tree_208;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_400 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_207),
 .b(tree_171),
 .c(tree_208)
);
wire [0:0] tree_209;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_401 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[10]),
 .b(in[176]),
 .c(tree_209)
);
wire [0:0] tree_210;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_402 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[31]),
 .b(in[191]),
 .c(tree_210)
);
wire [0:0] tree_211;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_403 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[11]),
 .b(in[167]),
 .c(tree_211)
);
wire [0:0] tree_212;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_404 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[50]),
 .b(in[143]),
 .c(tree_212)
);
wire [0:0] tree_213;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_405 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[86]),
 .b(1'h0),
 .c(tree_213)
);
wire [0:0] tree_214;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_406 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_213),
 .b(tree_138),
 .c(tree_214)
);
wire [0:0] tree_215;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_407 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[132]),
 .b(in[176]),
 .c(tree_215)
);
wire [0:0] tree_216;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_408 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[2]),
 .b(1'h0),
 .c(tree_216)
);
wire [0:0] tree_217;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_409 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_216),
 .b(tree_77),
 .c(tree_217)
);
wire [0:0] tree_218;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_410 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[43]),
 .b(in[174]),
 .c(tree_218)
);
wire [0:0] tree_219;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_411 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[106]),
 .b(1'h0),
 .c(tree_219)
);
wire [0:0] tree_220;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_412 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_219),
 .b(tree_89),
 .c(tree_220)
);
wire [0:0] tree_221;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_413 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[56]),
 .b(in[121]),
 .c(tree_221)
);
wire [0:0] tree_222;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_414 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[57]),
 .b(in[118]),
 .c(tree_222)
);
wire [0:0] tree_223;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_415 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[89]),
 .b(1'h0),
 .c(tree_223)
);
wire [0:0] tree_224;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_416 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_223),
 .b(tree_76),
 .c(tree_224)
);
wire [0:0] tree_225;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_417 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[16]),
 .b(in[53]),
 .c(tree_225)
);
wire [0:0] tree_226;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_418 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[129]),
 .b(in[158]),
 .c(tree_226)
);
wire [0:0] tree_227;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_419 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[81]),
 .b(in[139]),
 .c(tree_227)
);
wire [0:0] tree_228;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_420 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[94]),
 .b(in[182]),
 .c(tree_228)
);
wire [0:0] tree_229;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_421 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[78]),
 .b(1'h0),
 .c(tree_229)
);
wire [0:0] tree_230;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_422 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_229),
 .b(tree_10),
 .c(tree_230)
);
wire [0:0] tree_231;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_423 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[44]),
 .b(in[125]),
 .c(tree_231)
);
wire [0:0] tree_232;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_424 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[3]),
 .b(1'h0),
 .c(tree_232)
);
wire [0:0] tree_233;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_425 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_232),
 .b(tree_170),
 .c(tree_233)
);
wire [0:0] tree_234;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_426 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[58]),
 .b(in[154]),
 .c(tree_234)
);
wire [0:0] tree_235;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_427 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[25]),
 .b(in[27]),
 .c(tree_235)
);
wire [0:0] tree_236;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_428 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[107]),
 .b(in[147]),
 .c(tree_236)
);
wire [0:0] tree_237;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_429 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[160]),
 .b(in[162]),
 .c(tree_237)
);
wire [0:0] tree_238;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_430 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_205),
 .b(tree_70),
 .c(tree_238)
);
wire [0:0] tree_239;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_431 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[12]),
 .b(in[132]),
 .c(tree_239)
);
wire [0:0] tree_240;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_432 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[52]),
 .b(in[130]),
 .c(tree_240)
);
wire [0:0] tree_241;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_433 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[72]),
 .b(in[189]),
 .c(tree_241)
);
wire [0:0] tree_242;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_434 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[122]),
 .b(1'h0),
 .c(tree_242)
);
wire [0:0] tree_243;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_435 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_242),
 .b(tree_122),
 .c(tree_243)
);
wire [0:0] tree_244;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_436 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[145]),
 .b(in[187]),
 .c(tree_244)
);
wire [0:0] tree_245;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_437 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[26]),
 .b(in[28]),
 .c(tree_245)
);
wire [0:0] tree_246;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_438 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_7),
 .b(tree_227),
 .c(tree_246)
);
wire [0:0] tree_247;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_439 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[103]),
 .b(in[179]),
 .c(tree_247)
);
wire [0:0] tree_248;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_440 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[67]),
 .b(in[134]),
 .c(tree_248)
);
wire [0:0] tree_249;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_441 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[6]),
 .b(in[53]),
 .c(tree_249)
);
wire [0:0] tree_250;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_442 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[54]),
 .b(in[144]),
 .c(tree_250)
);
wire [0:0] tree_251;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_443 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[139]),
 .b(in[165]),
 .c(tree_251)
);
wire [0:0] tree_252;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_444 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[141]),
 .b(in[145]),
 .c(tree_252)
);
wire [0:0] tree_253;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_445 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[98]),
 .b(in[151]),
 .c(tree_253)
);
wire [0:0] tree_254;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_446 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[146]),
 .b(1'h0),
 .c(tree_254)
);
wire [0:0] tree_255;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_447 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_254),
 .b(tree_72),
 .c(tree_255)
);
wire [0:0] tree_256;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_448 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[15]),
 .b(1'h0),
 .c(tree_256)
);
wire [0:0] tree_257;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_449 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_256),
 .b(tree_60),
 .c(tree_257)
);
wire [0:0] tree_258;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_450 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[17]),
 .b(in[190]),
 .c(tree_258)
);
wire [0:0] tree_259;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_451 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[62]),
 .b(in[88]),
 .c(tree_259)
);
wire [0:0] tree_260;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_452 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[14]),
 .b(in[111]),
 .c(tree_260)
);
wire [0:0] tree_261;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_453 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[140]),
 .b(1'h0),
 .c(tree_261)
);
wire [0:0] tree_262;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_454 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_261),
 .b(tree_191),
 .c(tree_262)
);
wire [0:0] tree_263;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_455 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[155]),
 .b(in[168]),
 .c(tree_263)
);
wire [0:0] tree_264;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_456 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[31]),
 .b(in[156]),
 .c(tree_264)
);
wire [0:0] tree_265;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_457 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[38]),
 .b(in[161]),
 .c(tree_265)
);
wire [0:0] tree_266;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_458 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[113]),
 .b(in[126]),
 .c(tree_266)
);
wire [0:0] tree_267;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_459 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[80]),
 .b(1'h0),
 .c(tree_267)
);
wire [0:0] tree_268;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_460 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_267),
 .b(tree_86),
 .c(tree_268)
);
wire [0:0] tree_269;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_461 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[90]),
 .b(in[100]),
 .c(tree_269)
);
wire [0:0] tree_270;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_462 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[40]),
 .b(in[110]),
 .c(tree_270)
);
wire [0:0] tree_271;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_463 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[115]),
 .b(in[183]),
 .c(tree_271)
);
wire [0:0] tree_272;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_464 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[59]),
 .b(1'h0),
 .c(tree_272)
);
wire [0:0] tree_273;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_465 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_272),
 .b(tree_226),
 .c(tree_273)
);
wire [0:0] tree_274;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_466 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[20]),
 .b(in[98]),
 .c(tree_274)
);
wire [0:0] tree_275;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_467 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[114]),
 .b(in[155]),
 .c(tree_275)
);
wire [0:0] tree_276;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_468 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1),
 .b(tree_24),
 .c(tree_276)
);
wire [0:0] tree_277;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_469 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[9]),
 .b(in[75]),
 .c(tree_277)
);
wire [0:0] tree_278;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_470 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[63]),
 .b(in[161]),
 .c(tree_278)
);
wire [0:0] tree_279;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_471 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[48]),
 .b(in[148]),
 .c(tree_279)
);
wire [0:0] tree_280;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_472 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[69]),
 .b(in[187]),
 .c(tree_280)
);
wire [0:0] tree_281;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_473 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[138]),
 .b(in[190]),
 .c(tree_281)
);
wire [0:0] tree_282;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_474 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[64]),
 .b(in[145]),
 .c(tree_282)
);
wire [0:0] tree_283;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_475 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[38]),
 .b(1'h0),
 .c(tree_283)
);
wire [0:0] tree_284;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_476 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_283),
 .b(tree_38),
 .c(tree_284)
);
wire [0:0] tree_285;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_477 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[82]),
 .b(in[136]),
 .c(tree_285)
);
wire [0:0] tree_286;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_478 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[0]),
 .b(1'h0),
 .c(tree_286)
);
wire [0:0] tree_287;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_479 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_286),
 .b(tree_266),
 .c(tree_287)
);
wire [0:0] tree_288;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_480 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[14]),
 .b(1'h0),
 .c(tree_288)
);
wire [0:0] tree_289;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_481 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_288),
 .b(tree_201),
 .c(tree_289)
);
wire [0:0] tree_290;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_482 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[73]),
 .b(1'h0),
 .c(tree_290)
);
wire [0:0] tree_291;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_483 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_290),
 .b(tree_82),
 .c(tree_291)
);
wire [0:0] tree_292;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_484 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[97]),
 .b(in[150]),
 .c(tree_292)
);
wire [0:0] tree_293;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_485 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[28]),
 .b(1'h0),
 .c(tree_293)
);
wire [0:0] tree_294;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_486 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_293),
 .b(tree_73),
 .c(tree_294)
);
wire [0:0] tree_295;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_487 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[2]),
 .b(1'h0),
 .c(tree_295)
);
wire [0:0] tree_296;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_488 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_295),
 .b(tree_54),
 .c(tree_296)
);
wire [0:0] tree_297;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_489 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[43]),
 .b(1'h0),
 .c(tree_297)
);
wire [0:0] tree_298;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_490 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_297),
 .b(tree_194),
 .c(tree_298)
);
wire [0:0] tree_299;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_491 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[42]),
 .b(in[57]),
 .c(tree_299)
);
wire [0:0] tree_300;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_492 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[66]),
 .b(1'h0),
 .c(tree_300)
);
wire [0:0] tree_301;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_493 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_300),
 .b(tree_69),
 .c(tree_301)
);
wire [0:0] tree_302;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_494 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[20]),
 .b(in[45]),
 .c(tree_302)
);
wire [0:0] tree_303;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_495 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[140]),
 .b(1'h0),
 .c(tree_303)
);
wire [0:0] tree_304;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_496 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_303),
 .b(tree_165),
 .c(tree_304)
);
wire [0:0] tree_305;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_497 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[71]),
 .b(in[110]),
 .c(tree_305)
);
wire [0:0] tree_306;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_498 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[163]),
 .b(1'h0),
 .c(tree_306)
);
wire [0:0] tree_307;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_499 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_306),
 .b(tree_158),
 .c(tree_307)
);
wire [0:0] tree_308;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_500 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[189]),
 .b(1'h0),
 .c(tree_308)
);
wire [0:0] tree_309;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_501 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_308),
 .b(tree_28),
 .c(tree_309)
);
wire [0:0] tree_310;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_502 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[1]),
 .b(in[25]),
 .c(tree_310)
);
wire [0:0] tree_311;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_503 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[13]),
 .b(in[154]),
 .c(tree_311)
);
wire [0:0] tree_312;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_504 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[9]),
 .b(in[180]),
 .c(tree_312)
);
wire [0:0] tree_313;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_505 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[37]),
 .b(in[70]),
 .c(tree_313)
);
wire [0:0] tree_314;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_506 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[162]),
 .b(1'h0),
 .c(tree_314)
);
wire [0:0] tree_315;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_507 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_314),
 .b(tree_184),
 .c(tree_315)
);
wire [0:0] tree_316;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_508 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_46),
 .b(tree_274),
 .c(tree_316)
);
wire [0:0] tree_317;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_509 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[44]),
 .b(1'h0),
 .c(tree_317)
);
wire [0:0] tree_318;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_510 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_317),
 .b(tree_264),
 .c(tree_318)
);
wire [0:0] tree_319;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_511 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[33]),
 .b(in[128]),
 .c(tree_319)
);
wire [0:0] tree_320;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_512 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[79]),
 .b(in[125]),
 .c(tree_320)
);
wire [0:0] tree_321;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_513 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[117]),
 .b(in[120]),
 .c(tree_321)
);
wire [0:0] tree_322;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_514 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[62]),
 .b(in[130]),
 .c(tree_322)
);
wire [0:0] tree_323;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_515 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[132]),
 .b(in[186]),
 .c(tree_323)
);
wire [0:0] tree_324;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_516 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[189]),
 .b(1'h0),
 .c(tree_324)
);
wire [0:0] tree_325;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_517 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_324),
 .b(tree_3),
 .c(tree_325)
);
wire [0:0] tree_326;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_518 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[130]),
 .b(in[131]),
 .c(tree_326)
);
wire [0:0] tree_327;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_519 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[32]),
 .b(in[72]),
 .c(tree_327)
);
wire [0:0] tree_328;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_520 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[133]),
 .b(1'h0),
 .c(tree_328)
);
wire [0:0] tree_329;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_521 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_328),
 .b(tree_28),
 .c(tree_329)
);
wire [0:0] tree_330;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_522 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[31]),
 .b(in[34]),
 .c(tree_330)
);
wire [0:0] tree_331;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_523 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[92]),
 .b(in[157]),
 .c(tree_331)
);
wire [0:0] tree_332;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_524 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_159),
 .b(1'h0),
 .c(tree_332)
);
wire [0:0] tree_333;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_525 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_332),
 .b(tree_128),
 .c(tree_333)
);
wire [0:0] tree_334;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_526 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[116]),
 .b(in[117]),
 .c(tree_334)
);
wire [0:0] tree_335;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_527 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[127]),
 .b(in[167]),
 .c(tree_335)
);
wire [0:0] tree_336;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_528 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[7]),
 .b(in[76]),
 .c(tree_336)
);
wire [0:0] tree_337;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_529 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[6]),
 .b(in[58]),
 .c(tree_337)
);
wire [0:0] tree_338;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_530 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[31]),
 .b(in[108]),
 .c(tree_338)
);
wire [0:0] tree_339;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_531 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[34]),
 .b(in[186]),
 .c(tree_339)
);
wire [0:0] tree_340;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_532 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[178]),
 .b(1'h0),
 .c(tree_340)
);
wire [0:0] tree_341;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_533 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_340),
 .b(tree_172),
 .c(tree_341)
);
wire [0:0] tree_342;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_534 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[12]),
 .b(in[50]),
 .c(tree_342)
);
wire [0:0] tree_343;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_535 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[13]),
 .b(1'h0),
 .c(tree_343)
);
wire [0:0] tree_344;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_536 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_343),
 .b(tree_103),
 .c(tree_344)
);
wire [0:0] tree_345;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_537 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[2]),
 .b(1'h0),
 .c(tree_345)
);
wire [0:0] tree_346;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_538 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_345),
 .b(tree_245),
 .c(tree_346)
);
wire [0:0] tree_347;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_539 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[32]),
 .b(in[122]),
 .c(tree_347)
);
wire [0:0] tree_348;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_540 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_88),
 .b(1'h0),
 .c(tree_348)
);
wire [0:0] tree_349;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_541 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_348),
 .b(tree_208),
 .c(tree_349)
);
wire [0:0] tree_350;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_542 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[74]),
 .b(1'h0),
 .c(tree_350)
);
wire [0:0] tree_351;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_543 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_350),
 .b(tree_152),
 .c(tree_351)
);
wire [0:0] tree_352;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_544 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[85]),
 .b(1'h0),
 .c(tree_352)
);
wire [0:0] tree_353;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_545 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_352),
 .b(tree_86),
 .c(tree_353)
);
wire [0:0] tree_354;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_546 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[108]),
 .b(in[128]),
 .c(tree_354)
);
wire [0:0] tree_355;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_547 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[4]),
 .b(in[177]),
 .c(tree_355)
);
wire [0:0] tree_356;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_548 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[82]),
 .b(in[110]),
 .c(tree_356)
);
wire [0:0] tree_357;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_549 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_43),
 .b(tree_335),
 .c(tree_357)
);
wire [0:0] tree_358;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_550 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[56]),
 .b(in[150]),
 .c(tree_358)
);
wire [0:0] tree_359;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_551 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[29]),
 .b(in[151]),
 .c(tree_359)
);
wire [0:0] tree_360;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_552 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[44]),
 .b(in[59]),
 .c(tree_360)
);
wire [0:0] tree_361;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_553 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[47]),
 .b(in[156]),
 .c(tree_361)
);
wire [0:0] tree_362;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_554 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[92]),
 .b(in[106]),
 .c(tree_362)
);
wire [0:0] tree_363;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_555 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[88]),
 .b(1'h0),
 .c(tree_363)
);
wire [0:0] tree_364;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_556 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_363),
 .b(tree_68),
 .c(tree_364)
);
wire [0:0] tree_365;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_557 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_105),
 .b(tree_311),
 .c(tree_365)
);
wire [0:0] tree_366;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_558 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[96]),
 .b(in[137]),
 .c(tree_366)
);
wire [0:0] tree_367;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_559 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[10]),
 .b(in[75]),
 .c(tree_367)
);
wire [0:0] tree_368;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_560 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[70]),
 .b(in[79]),
 .c(tree_368)
);
wire [0:0] tree_369;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_561 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[156]),
 .b(1'h0),
 .c(tree_369)
);
wire [0:0] tree_370;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_562 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_369),
 .b(tree_327),
 .c(tree_370)
);
wire [0:0] tree_371;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_563 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[174]),
 .b(1'h0),
 .c(tree_371)
);
wire [0:0] tree_372;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_564 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_371),
 .b(tree_33),
 .c(tree_372)
);
wire [0:0] tree_373;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_565 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[15]),
 .b(1'h0),
 .c(tree_373)
);
wire [0:0] tree_374;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_566 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_373),
 .b(1'h0),
 .c(tree_374)
);
wire [0:0] tree_375;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_567 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_374),
 .b(tree_344),
 .c(tree_375)
);
wire [0:0] tree_376;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_568 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[1]),
 .b(in[136]),
 .c(tree_376)
);
wire [0:0] tree_377;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_569 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[159]),
 .b(in[169]),
 .c(tree_377)
);
wire [0:0] tree_378;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_570 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[131]),
 .b(in[163]),
 .c(tree_378)
);
wire [0:0] tree_379;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_571 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[5]),
 .b(in[123]),
 .c(tree_379)
);
wire [0:0] tree_380;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_572 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[177]),
 .b(in[181]),
 .c(tree_380)
);
wire [0:0] tree_381;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_573 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[148]),
 .b(1'h0),
 .c(tree_381)
);
wire [0:0] tree_382;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_574 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_381),
 .b(tree_336),
 .c(tree_382)
);
wire [0:0] tree_383;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_575 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[149]),
 .b(in[178]),
 .c(tree_383)
);
wire [0:0] tree_384;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_576 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[187]),
 .b(1'h0),
 .c(tree_384)
);
wire [0:0] tree_385;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_577 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_384),
 .b(tree_151),
 .c(tree_385)
);
wire [0:0] tree_386;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_578 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[119]),
 .b(in[126]),
 .c(tree_386)
);
wire [0:0] tree_387;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_579 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[55]),
 .b(in[82]),
 .c(tree_387)
);
wire [0:0] tree_388;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_580 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[77]),
 .b(1'h0),
 .c(tree_388)
);
wire [0:0] tree_389;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_581 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_388),
 .b(tree_15),
 .c(tree_389)
);
wire [0:0] tree_390;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_582 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[138]),
 .b(1'h0),
 .c(tree_390)
);
wire [0:0] tree_391;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_583 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_390),
 .b(tree_108),
 .c(tree_391)
);
wire [0:0] tree_392;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_584 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[50]),
 .b(in[174]),
 .c(tree_392)
);
wire [0:0] tree_393;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_585 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[62]),
 .b(1'h0),
 .c(tree_393)
);
wire [0:0] tree_394;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_586 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_393),
 .b(tree_79),
 .c(tree_394)
);
wire [0:0] tree_395;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_587 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[16]),
 .b(in[137]),
 .c(tree_395)
);
wire [0:0] tree_396;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_588 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[95]),
 .b(in[188]),
 .c(tree_396)
);
wire [0:0] tree_397;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_589 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[53]),
 .b(in[84]),
 .c(tree_397)
);
wire [0:0] tree_398;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_590 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[46]),
 .b(1'h0),
 .c(tree_398)
);
wire [0:0] tree_399;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_591 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_398),
 .b(tree_190),
 .c(tree_399)
);
wire [0:0] tree_400;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_592 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[40]),
 .b(in[124]),
 .c(tree_400)
);
wire [0:0] tree_401;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_593 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[21]),
 .b(in[35]),
 .c(tree_401)
);
wire [0:0] tree_402;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_594 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[59]),
 .b(in[166]),
 .c(tree_402)
);
wire [0:0] tree_403;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_595 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[77]),
 .b(in[144]),
 .c(tree_403)
);
wire [0:0] tree_404;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_596 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[117]),
 .b(in[141]),
 .c(tree_404)
);
wire [0:0] tree_405;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_597 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[159]),
 .b(in[189]),
 .c(tree_405)
);
wire [0:0] tree_406;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_598 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[11]),
 .b(in[105]),
 .c(tree_406)
);
wire [0:0] tree_407;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_599 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[38]),
 .b(1'h0),
 .c(tree_407)
);
wire [0:0] tree_408;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_600 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_407),
 .b(tree_29),
 .c(tree_408)
);
wire [0:0] tree_409;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_601 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[8]),
 .b(in[127]),
 .c(tree_409)
);
wire [0:0] tree_410;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_602 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[15]),
 .b(in[81]),
 .c(tree_410)
);
wire [0:0] tree_411;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_603 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_339),
 .b(tree_42),
 .c(tree_411)
);
wire [0:0] tree_412;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_604 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[55]),
 .b(in[148]),
 .c(tree_412)
);
wire [0:0] tree_413;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_605 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_10),
 .b(tree_263),
 .c(tree_413)
);
wire [0:0] tree_414;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_606 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[100]),
 .b(1'h0),
 .c(tree_414)
);
wire [0:0] tree_415;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_607 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_414),
 .b(tree_30),
 .c(tree_415)
);
wire [0:0] tree_416;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_608 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[76]),
 .b(in[166]),
 .c(tree_416)
);
wire [0:0] tree_417;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_609 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[56]),
 .b(1'h0),
 .c(tree_417)
);
wire [0:0] tree_418;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_610 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_417),
 .b(tree_205),
 .c(tree_418)
);
wire [0:0] tree_419;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_611 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[58]),
 .b(1'h0),
 .c(tree_419)
);
wire [0:0] tree_420;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_612 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_419),
 .b(tree_88),
 .c(tree_420)
);
wire [0:0] tree_421;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_613 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[134]),
 .b(1'h0),
 .c(tree_421)
);
wire [0:0] tree_422;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_614 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_421),
 .b(tree_0),
 .c(tree_422)
);
wire [0:0] tree_423;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_615 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_106),
 .b(tree_331),
 .c(tree_423)
);
wire [0:0] tree_424;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_616 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[1]),
 .b(1'h0),
 .c(tree_424)
);
wire [0:0] tree_425;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_617 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_424),
 .b(tree_68),
 .c(tree_425)
);
wire [0:0] tree_426;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_618 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[61]),
 .b(in[83]),
 .c(tree_426)
);
wire [0:0] tree_427;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_619 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[67]),
 .b(1'h0),
 .c(tree_427)
);
wire [0:0] tree_428;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_620 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_427),
 .b(tree_32),
 .c(tree_428)
);
wire [0:0] tree_429;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_621 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_327),
 .b(tree_251),
 .c(tree_429)
);
wire [0:0] tree_430;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_622 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_46),
 .b(tree_97),
 .c(tree_430)
);
wire [0:0] tree_431;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_623 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_3),
 .b(tree_102),
 .c(tree_431)
);
wire [0:0] tree_432;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_624 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_181),
 .b(tree_183),
 .c(tree_432)
);
wire [0:0] tree_433;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_625 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[10]),
 .b(1'h0),
 .c(tree_433)
);
wire [0:0] tree_434;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_626 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_433),
 .b(tree_22),
 .c(tree_434)
);
wire [0:0] tree_435;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_627 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[185]),
 .b(1'h0),
 .c(tree_435)
);
wire [0:0] tree_436;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_628 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_435),
 .b(tree_96),
 .c(tree_436)
);
wire [0:0] tree_437;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_629 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[34]),
 .b(1'h0),
 .c(tree_437)
);
wire [0:0] tree_438;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_630 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_437),
 .b(tree_193),
 .c(tree_438)
);
wire [0:0] tree_439;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_631 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[111]),
 .b(1'h0),
 .c(tree_439)
);
wire [0:0] tree_440;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_632 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_439),
 .b(tree_16),
 .c(tree_440)
);
wire [0:0] tree_441;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_633 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[137]),
 .b(1'h0),
 .c(tree_441)
);
wire [0:0] tree_442;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_634 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_441),
 .b(tree_91),
 .c(tree_442)
);
wire [0:0] tree_443;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_635 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[157]),
 .b(1'h0),
 .c(tree_443)
);
wire [0:0] tree_444;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_636 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_443),
 .b(tree_106),
 .c(tree_444)
);
wire [0:0] tree_445;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_637 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[18]),
 .b(in[186]),
 .c(tree_445)
);
wire [0:0] tree_446;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_638 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_50),
 .b(1'h0),
 .c(tree_446)
);
wire [0:0] tree_447;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_639 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_446),
 .b(tree_408),
 .c(tree_447)
);
wire [0:0] tree_448;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_640 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[169]),
 .b(in[184]),
 .c(tree_448)
);
wire [0:0] tree_449;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_641 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[152]),
 .b(1'h0),
 .c(tree_449)
);
wire [0:0] tree_450;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_642 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_449),
 .b(tree_151),
 .c(tree_450)
);
wire [0:0] tree_451;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_643 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[57]),
 .b(1'h0),
 .c(tree_451)
);
wire [0:0] tree_452;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_644 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_451),
 .b(tree_360),
 .c(tree_452)
);
wire [0:0] tree_453;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_645 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[102]),
 .b(in[106]),
 .c(tree_453)
);
wire [0:0] tree_454;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_646 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[22]),
 .b(1'h0),
 .c(tree_454)
);
wire [0:0] tree_455;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_647 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_454),
 .b(1'h0),
 .c(tree_455)
);
wire [0:0] tree_456;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_648 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_455),
 .b(tree_434),
 .c(tree_456)
);
wire [0:0] tree_457;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_649 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[35]),
 .b(in[153]),
 .c(tree_457)
);
wire [0:0] tree_458;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_650 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[51]),
 .b(1'h0),
 .c(tree_458)
);
wire [0:0] tree_459;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_651 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_458),
 .b(tree_61),
 .c(tree_459)
);
wire [0:0] tree_460;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_652 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[33]),
 .b(in[41]),
 .c(tree_460)
);
wire [0:0] tree_461;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_653 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[47]),
 .b(in[73]),
 .c(tree_461)
);
wire [0:0] tree_462;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_654 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[98]),
 .b(in[136]),
 .c(tree_462)
);
wire [0:0] tree_463;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_655 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[28]),
 .b(in[166]),
 .c(tree_463)
);
wire [0:0] tree_464;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_656 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_358),
 .b(tree_448),
 .c(tree_464)
);
wire [0:0] tree_465;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_657 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[14]),
 .b(in[96]),
 .c(tree_465)
);
wire [0:0] tree_466;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_658 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[87]),
 .b(1'h0),
 .c(tree_466)
);
wire [0:0] tree_467;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_659 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_466),
 .b(tree_281),
 .c(tree_467)
);
wire [0:0] tree_468;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_660 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[155]),
 .b(1'h0),
 .c(tree_468)
);
wire [0:0] tree_469;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_661 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_468),
 .b(tree_163),
 .c(tree_469)
);
wire [0:0] tree_470;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_662 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[51]),
 .b(in[174]),
 .c(tree_470)
);
wire [0:0] tree_471;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_663 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[68]),
 .b(in[123]),
 .c(tree_471)
);
wire [0:0] tree_472;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_664 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[113]),
 .b(1'h0),
 .c(tree_472)
);
wire [0:0] tree_473;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_665 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_472),
 .b(tree_277),
 .c(tree_473)
);
wire [0:0] tree_474;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_666 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[185]),
 .b(1'h0),
 .c(tree_474)
);
wire [0:0] tree_475;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_667 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_474),
 .b(tree_198),
 .c(tree_475)
);
wire [0:0] tree_476;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_668 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[124]),
 .b(in[172]),
 .c(tree_476)
);
wire [0:0] tree_477;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_669 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[151]),
 .b(1'h0),
 .c(tree_477)
);
wire [0:0] tree_478;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_670 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_477),
 .b(tree_247),
 .c(tree_478)
);
wire [0:0] tree_479;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_671 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[175]),
 .b(1'h0),
 .c(tree_479)
);
wire [0:0] tree_480;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_672 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_479),
 .b(tree_43),
 .c(tree_480)
);
wire [0:0] tree_481;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_673 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_465),
 .b(1'h0),
 .c(tree_481)
);
wire [0:0] tree_482;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_674 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_415),
 .b(tree_481),
 .c(tree_482)
);
wire [0:0] tree_483;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_675 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[26]),
 .b(in[182]),
 .c(tree_483)
);
wire [0:0] tree_484;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_676 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[6]),
 .b(1'h0),
 .c(tree_484)
);
wire [0:0] tree_485;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_677 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_484),
 .b(tree_76),
 .c(tree_485)
);
wire [0:0] tree_486;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_678 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[157]),
 .b(1'h0),
 .c(tree_486)
);
wire [0:0] tree_487;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_679 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_486),
 .b(tree_140),
 .c(tree_487)
);
wire [0:0] tree_488;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_680 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_99),
 .b(tree_201),
 .c(tree_488)
);
wire [0:0] tree_489;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_681 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[18]),
 .b(in[79]),
 .c(tree_489)
);
wire [0:0] tree_490;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_682 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[33]),
 .b(in[172]),
 .c(tree_490)
);
wire [0:0] tree_491;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_683 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[31]),
 .b(1'h0),
 .c(tree_491)
);
wire [0:0] tree_492;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_684 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_491),
 .b(tree_33),
 .c(tree_492)
);
wire [0:0] tree_493;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_685 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[37]),
 .b(1'h0),
 .c(tree_493)
);
wire [0:0] tree_494;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_686 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_493),
 .b(tree_48),
 .c(tree_494)
);
wire [0:0] tree_495;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_687 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[153]),
 .b(1'h0),
 .c(tree_495)
);
wire [0:0] tree_496;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_688 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_495),
 .b(tree_400),
 .c(tree_496)
);
wire [0:0] tree_497;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_689 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[179]),
 .b(1'h0),
 .c(tree_497)
);
wire [0:0] tree_498;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_690 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_497),
 .b(1'h0),
 .c(tree_498)
);
wire [0:0] tree_499;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_691 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_498),
 .b(tree_434),
 .c(tree_499)
);
wire [0:0] tree_500;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_692 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[90]),
 .b(1'h0),
 .c(tree_500)
);
wire [0:0] tree_501;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_693 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_500),
 .b(tree_189),
 .c(tree_501)
);
wire [0:0] tree_502;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_694 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[21]),
 .b(in[72]),
 .c(tree_502)
);
wire [0:0] tree_503;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_695 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[84]),
 .b(1'h0),
 .c(tree_503)
);
wire [0:0] tree_504;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_696 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_503),
 .b(tree_9),
 .c(tree_504)
);
wire [0:0] tree_505;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_697 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[60]),
 .b(1'h0),
 .c(tree_505)
);
wire [0:0] tree_506;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_698 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_505),
 .b(tree_305),
 .c(tree_506)
);
wire [0:0] tree_507;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_699 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_211),
 .b(tree_235),
 .c(tree_507)
);
wire [0:0] tree_508;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_700 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[73]),
 .b(in[88]),
 .c(tree_508)
);
wire [0:0] tree_509;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_701 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_26),
 .b(tree_470),
 .c(tree_509)
);
wire [0:0] tree_510;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_702 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[9]),
 .b(in[53]),
 .c(tree_510)
);
wire [0:0] tree_511;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_703 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_334),
 .b(tree_141),
 .c(tree_511)
);
wire [0:0] tree_512;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_704 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[0]),
 .b(1'h0),
 .c(tree_512)
);
wire [0:0] tree_513;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_705 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_512),
 .b(tree_80),
 .c(tree_513)
);
wire [0:0] tree_514;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_706 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[161]),
 .b(1'h0),
 .c(tree_514)
);
wire [0:0] tree_515;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_707 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_514),
 .b(tree_82),
 .c(tree_515)
);
wire [0:0] tree_516;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_708 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[181]),
 .b(1'h0),
 .c(tree_516)
);
wire [0:0] tree_517;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_709 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_516),
 .b(tree_299),
 .c(tree_517)
);
wire [0:0] tree_518;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_710 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[117]),
 .b(in[164]),
 .c(tree_518)
);
wire [0:0] tree_519;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_711 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_14),
 .b(tree_156),
 .c(tree_519)
);
wire [0:0] tree_520;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_712 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_277),
 .b(1'h0),
 .c(tree_520)
);
wire [0:0] tree_521;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_713 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_520),
 .b(tree_440),
 .c(tree_521)
);
wire [0:0] tree_522;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_714 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_106),
 .b(tree_383),
 .c(tree_522)
);
wire [0:0] tree_523;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_715 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[70]),
 .b(in[142]),
 .c(tree_523)
);
wire [0:0] tree_524;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_716 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[185]),
 .b(1'h0),
 .c(tree_524)
);
wire [0:0] tree_525;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_717 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_524),
 .b(tree_157),
 .c(tree_525)
);
wire [0:0] tree_526;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_718 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[93]),
 .b(in[96]),
 .c(tree_526)
);
wire [0:0] tree_527;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_719 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[4]),
 .b(1'h0),
 .c(tree_527)
);
wire [0:0] tree_528;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_720 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_527),
 .b(1'h0),
 .c(tree_528)
);
wire [0:0] tree_529;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_721 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_528),
 .b(tree_154),
 .c(tree_529)
);
wire [0:0] tree_530;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_722 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[17]),
 .b(1'h0),
 .c(tree_530)
);
wire [0:0] tree_531;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_723 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_530),
 .b(tree_190),
 .c(tree_531)
);
wire [0:0] tree_532;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_724 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[56]),
 .b(in[64]),
 .c(tree_532)
);
wire [0:0] tree_533;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_725 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[127]),
 .b(1'h0),
 .c(tree_533)
);
wire [0:0] tree_534;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_726 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_533),
 .b(tree_275),
 .c(tree_534)
);
wire [0:0] tree_535;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_727 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[136]),
 .b(1'h0),
 .c(tree_535)
);
wire [0:0] tree_536;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_728 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_535),
 .b(tree_168),
 .c(tree_536)
);
wire [0:0] tree_537;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_729 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[158]),
 .b(in[173]),
 .c(tree_537)
);
wire [0:0] tree_538;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_730 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_22),
 .b(1'h0),
 .c(tree_538)
);
wire [0:0] tree_539;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_731 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_538),
 .b(tree_325),
 .c(tree_539)
);
wire [0:0] tree_540;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_732 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[186]),
 .b(1'h0),
 .c(tree_540)
);
wire [0:0] tree_541;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_733 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_540),
 .b(tree_274),
 .c(tree_541)
);
wire [0:0] tree_542;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_734 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[24]),
 .b(in[133]),
 .c(tree_542)
);
wire [0:0] tree_543;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_735 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_165),
 .b(tree_188),
 .c(tree_543)
);
wire [0:0] tree_544;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_736 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[7]),
 .b(in[113]),
 .c(tree_544)
);
wire [0:0] tree_545;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_737 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[11]),
 .b(1'h0),
 .c(tree_545)
);
wire [0:0] tree_546;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_738 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_545),
 .b(tree_25),
 .c(tree_546)
);
wire [0:0] tree_547;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_739 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[68]),
 .b(in[85]),
 .c(tree_547)
);
wire [0:0] tree_548;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_740 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[111]),
 .b(1'h0),
 .c(tree_548)
);
wire [0:0] tree_549;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_741 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_548),
 .b(tree_87),
 .c(tree_549)
);
wire [0:0] tree_550;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_742 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[3]),
 .b(in[24]),
 .c(tree_550)
);
wire [0:0] tree_551;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_743 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[65]),
 .b(1'h0),
 .c(tree_551)
);
wire [0:0] tree_552;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_744 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_551),
 .b(tree_100),
 .c(tree_552)
);
wire [0:0] tree_553;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_745 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[183]),
 .b(1'h0),
 .c(tree_553)
);
wire [0:0] tree_554;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_746 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_553),
 .b(tree_7),
 .c(tree_554)
);
wire [0:0] tree_555;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_747 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_122),
 .b(1'h0),
 .c(tree_555)
);
wire [0:0] tree_556;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_748 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_555),
 .b(tree_175),
 .c(tree_556)
);
wire [0:0] tree_557;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_749 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[92]),
 .b(1'h0),
 .c(tree_557)
);
wire [0:0] tree_558;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_750 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_557),
 .b(tree_107),
 .c(tree_558)
);
wire [0:0] tree_559;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_751 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[83]),
 .b(in[165]),
 .c(tree_559)
);
wire [0:0] tree_560;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_752 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_104),
 .b(tree_71),
 .c(tree_560)
);
wire [0:0] tree_561;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_753 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[167]),
 .b(1'h0),
 .c(tree_561)
);
wire [0:0] tree_562;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_754 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_561),
 .b(tree_14),
 .c(tree_562)
);
wire [0:0] tree_563;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_755 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_285),
 .b(tree_0),
 .c(tree_563)
);
wire [0:0] tree_564;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_756 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[12]),
 .b(1'h0),
 .c(tree_564)
);
wire [0:0] tree_565;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_757 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_564),
 .b(tree_383),
 .c(tree_565)
);
wire [0:0] tree_566;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_758 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[54]),
 .b(in[66]),
 .c(tree_566)
);
wire [0:0] tree_567;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_759 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[99]),
 .b(1'h0),
 .c(tree_567)
);
wire [0:0] tree_568;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_760 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_567),
 .b(1'h0),
 .c(tree_568)
);
wire [0:0] tree_569;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_761 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_568),
 .b(tree_95),
 .c(tree_569)
);
wire [0:0] tree_570;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_762 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[173]),
 .b(1'h0),
 .c(tree_570)
);
wire [0:0] tree_571;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_763 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_570),
 .b(tree_137),
 .c(tree_571)
);
wire [0:0] tree_572;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_764 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[8]),
 .b(in[190]),
 .c(tree_572)
);
wire [0:0] tree_573;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_765 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[151]),
 .b(1'h0),
 .c(tree_573)
);
wire [0:0] tree_574;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_766 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_573),
 .b(tree_7),
 .c(tree_574)
);
wire [0:0] tree_575;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_767 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[42]),
 .b(1'h0),
 .c(tree_575)
);
wire [0:0] tree_576;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_768 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_575),
 .b(tree_160),
 .c(tree_576)
);
wire [0:0] tree_577;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_769 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[89]),
 .b(in[116]),
 .c(tree_577)
);
wire [0:0] tree_578;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_770 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_360),
 .b(tree_194),
 .c(tree_578)
);
wire [0:0] tree_579;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_771 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[23]),
 .b(in[127]),
 .c(tree_579)
);
wire [0:0] tree_580;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_772 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[9]),
 .b(in[22]),
 .c(tree_580)
);
wire [0:0] tree_581;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_773 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[85]),
 .b(1'h0),
 .c(tree_581)
);
wire [0:0] tree_582;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_774 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_581),
 .b(tree_205),
 .c(tree_582)
);
wire [0:0] tree_583;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_775 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[13]),
 .b(in[45]),
 .c(tree_583)
);
wire [0:0] tree_584;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_776 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_103),
 .b(tree_310),
 .c(tree_584)
);
wire [0:0] tree_585;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_777 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_165),
 .b(tree_323),
 .c(tree_585)
);
wire [0:0] tree_586;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_778 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[78]),
 .b(1'h0),
 .c(tree_586)
);
wire [0:0] tree_587;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_779 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_586),
 .b(tree_23),
 .c(tree_587)
);
wire [0:0] tree_588;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_780 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[81]),
 .b(in[142]),
 .c(tree_588)
);
wire [0:0] tree_589;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_781 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[61]),
 .b(1'h0),
 .c(tree_589)
);
wire [0:0] tree_590;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_782 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_589),
 .b(tree_13),
 .c(tree_590)
);
wire [0:0] tree_591;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_783 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_107),
 .b(tree_281),
 .c(tree_591)
);
wire [0:0] tree_592;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_784 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_266),
 .b(tree_401),
 .c(tree_592)
);
wire [0:0] tree_593;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_785 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[23]),
 .b(in[46]),
 .c(tree_593)
);
wire [0:0] tree_594;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_786 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[97]),
 .b(in[162]),
 .c(tree_594)
);
wire [0:0] tree_595;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_787 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_59),
 .b(tree_52),
 .c(tree_595)
);
wire [0:0] tree_596;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_788 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[0]),
 .b(in[157]),
 .c(tree_596)
);
wire [0:0] tree_597;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_789 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[91]),
 .b(1'h0),
 .c(tree_597)
);
wire [0:0] tree_598;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_790 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_597),
 .b(tree_339),
 .c(tree_598)
);
wire [0:0] tree_599;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_791 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[36]),
 .b(in[55]),
 .c(tree_599)
);
wire [0:0] tree_600;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_792 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_39),
 .b(tree_2),
 .c(tree_600)
);
wire [0:0] tree_601;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_793 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[7]),
 .b(in[99]),
 .c(tree_601)
);
wire [0:0] tree_602;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_794 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[134]),
 .b(in[176]),
 .c(tree_602)
);
wire [0:0] tree_603;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_795 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[95]),
 .b(in[107]),
 .c(tree_603)
);
wire [0:0] tree_604;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_796 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[54]),
 .b(1'h0),
 .c(tree_604)
);
wire [0:0] tree_605;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_797 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_604),
 .b(tree_50),
 .c(tree_605)
);
wire [0:0] tree_606;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_798 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[72]),
 .b(in[114]),
 .c(tree_606)
);
wire [0:0] tree_607;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_799 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[129]),
 .b(1'h0),
 .c(tree_607)
);
wire [0:0] tree_608;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_800 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_607),
 .b(tree_180),
 .c(tree_608)
);
wire [0:0] tree_609;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_801 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_526),
 .b(tree_17),
 .c(tree_609)
);
wire [0:0] tree_610;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_802 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_173),
 .b(tree_51),
 .c(tree_610)
);
wire [0:0] tree_611;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_803 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[100]),
 .b(1'h0),
 .c(tree_611)
);
wire [0:0] tree_612;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_804 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_611),
 .b(tree_4),
 .c(tree_612)
);
wire [0:0] tree_613;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_805 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_137),
 .b(tree_577),
 .c(tree_613)
);
wire [0:0] tree_614;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_806 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[24]),
 .b(in[127]),
 .c(tree_614)
);
wire [0:0] tree_615;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_807 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[112]),
 .b(1'h0),
 .c(tree_615)
);
wire [0:0] tree_616;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_808 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_615),
 .b(tree_104),
 .c(tree_616)
);
wire [0:0] tree_617;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_809 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[165]),
 .b(1'h0),
 .c(tree_617)
);
wire [0:0] tree_618;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_810 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_617),
 .b(tree_376),
 .c(tree_618)
);
wire [0:0] tree_619;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_811 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[94]),
 .b(1'h0),
 .c(tree_619)
);
wire [0:0] tree_620;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_812 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_619),
 .b(tree_44),
 .c(tree_620)
);
wire [0:0] tree_621;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_813 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[123]),
 .b(in[191]),
 .c(tree_621)
);
wire [0:0] tree_622;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_814 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[22]),
 .b(in[177]),
 .c(tree_622)
);
wire [0:0] tree_623;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_815 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[130]),
 .b(1'h0),
 .c(tree_623)
);
wire [0:0] tree_624;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_816 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_623),
 .b(tree_211),
 .c(tree_624)
);
wire [0:0] tree_625;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_817 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_164),
 .b(1'h0),
 .c(tree_625)
);
wire [0:0] tree_626;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_818 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_625),
 .b(tree_576),
 .c(tree_626)
);
wire [0:0] tree_627;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_819 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[32]),
 .b(1'h0),
 .c(tree_627)
);
wire [0:0] tree_628;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_820 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_627),
 .b(tree_22),
 .c(tree_628)
);
wire [0:0] tree_629;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_821 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_0),
 .b(tree_132),
 .c(tree_629)
);
wire [0:0] tree_630;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_822 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[159]),
 .b(1'h0),
 .c(tree_630)
);
wire [0:0] tree_631;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_823 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_630),
 .b(tree_156),
 .c(tree_631)
);
wire [0:0] tree_632;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_824 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[6]),
 .b(in[79]),
 .c(tree_632)
);
wire [0:0] tree_633;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_825 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_83),
 .b(tree_326),
 .c(tree_633)
);
wire [0:0] tree_634;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_826 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[48]),
 .b(in[55]),
 .c(tree_634)
);
wire [0:0] tree_635;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_827 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[141]),
 .b(1'h0),
 .c(tree_635)
);
wire [0:0] tree_636;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_828 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_635),
 .b(tree_70),
 .c(tree_636)
);
wire [0:0] tree_637;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_829 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[145]),
 .b(1'h0),
 .c(tree_637)
);
wire [0:0] tree_638;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_830 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_637),
 .b(tree_583),
 .c(tree_638)
);
wire [0:0] tree_639;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_831 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[168]),
 .b(1'h0),
 .c(tree_639)
);
wire [0:0] tree_640;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_832 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_639),
 .b(1'h0),
 .c(tree_640)
);
wire [0:0] tree_641;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_833 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_640),
 .b(tree_214),
 .c(tree_641)
);
wire [0:0] tree_642;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_834 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_305),
 .b(1'h0),
 .c(tree_642)
);
wire [0:0] tree_643;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_835 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_642),
 .b(tree_475),
 .c(tree_643)
);
wire [0:0] tree_644;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_836 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[61]),
 .b(1'h0),
 .c(tree_644)
);
wire [0:0] tree_645;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_837 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_644),
 .b(tree_234),
 .c(tree_645)
);
wire [0:0] tree_646;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_838 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_205),
 .b(tree_137),
 .c(tree_646)
);
wire [0:0] tree_647;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_839 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[152]),
 .b(1'h0),
 .c(tree_647)
);
wire [0:0] tree_648;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_840 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_647),
 .b(tree_14),
 .c(tree_648)
);
wire [0:0] tree_649;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_841 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_15),
 .b(tree_81),
 .c(tree_649)
);
wire [0:0] tree_650;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_842 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[46]),
 .b(1'h0),
 .c(tree_650)
);
wire [0:0] tree_651;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_843 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_650),
 .b(tree_9),
 .c(tree_651)
);
wire [0:0] tree_652;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_844 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[49]),
 .b(in[103]),
 .c(tree_652)
);
wire [0:0] tree_653;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_845 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[68]),
 .b(in[145]),
 .c(tree_653)
);
wire [0:0] tree_654;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_846 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[59]),
 .b(1'h0),
 .c(tree_654)
);
wire [0:0] tree_655;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_847 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_654),
 .b(tree_270),
 .c(tree_655)
);
wire [0:0] tree_656;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_848 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_153),
 .b(tree_250),
 .c(tree_656)
);
wire [0:0] tree_657;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_849 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[19]),
 .b(1'h0),
 .c(tree_657)
);
wire [0:0] tree_658;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_850 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_657),
 .b(tree_105),
 .c(tree_658)
);
wire [0:0] tree_659;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_851 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[119]),
 .b(1'h0),
 .c(tree_659)
);
wire [0:0] tree_660;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_852 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_659),
 .b(tree_281),
 .c(tree_660)
);
wire [0:0] tree_661;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_853 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_5),
 .b(tree_152),
 .c(tree_661)
);
wire [0:0] tree_662;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_854 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[71]),
 .b(1'h0),
 .c(tree_662)
);
wire [0:0] tree_663;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_855 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_662),
 .b(tree_173),
 .c(tree_663)
);
wire [0:0] tree_664;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_856 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[7]),
 .b(1'h0),
 .c(tree_664)
);
wire [0:0] tree_665;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_857 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_664),
 .b(tree_263),
 .c(tree_665)
);
wire [0:0] tree_666;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_858 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[179]),
 .b(1'h0),
 .c(tree_666)
);
wire [0:0] tree_667;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_859 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_666),
 .b(tree_34),
 .c(tree_667)
);
wire [0:0] tree_668;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_860 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_185),
 .b(tree_355),
 .c(tree_668)
);
wire [0:0] tree_669;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_861 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[0]),
 .b(1'h0),
 .c(tree_669)
);
wire [0:0] tree_670;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_862 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_669),
 .b(tree_89),
 .c(tree_670)
);
wire [0:0] tree_671;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_863 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[26]),
 .b(1'h0),
 .c(tree_671)
);
wire [0:0] tree_672;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_864 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_671),
 .b(tree_120),
 .c(tree_672)
);
wire [0:0] tree_673;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_865 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[186]),
 .b(1'h0),
 .c(tree_673)
);
wire [0:0] tree_674;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_866 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_673),
 .b(1'h0),
 .c(tree_674)
);
wire [0:0] tree_675;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_867 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_674),
 .b(tree_612),
 .c(tree_675)
);
wire [0:0] tree_676;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_868 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[75]),
 .b(1'h0),
 .c(tree_676)
);
wire [0:0] tree_677;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_869 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_676),
 .b(tree_101),
 .c(tree_677)
);
wire [0:0] tree_678;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_870 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[40]),
 .b(in[76]),
 .c(tree_678)
);
wire [0:0] tree_679;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_871 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[119]),
 .b(1'h0),
 .c(tree_679)
);
wire [0:0] tree_680;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_872 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_679),
 .b(tree_35),
 .c(tree_680)
);
wire [0:0] tree_681;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_873 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_38),
 .b(tree_180),
 .c(tree_681)
);
wire [0:0] tree_682;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_874 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[5]),
 .b(1'h0),
 .c(tree_682)
);
wire [0:0] tree_683;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_875 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_682),
 .b(tree_270),
 .c(tree_683)
);
wire [0:0] tree_684;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_876 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[42]),
 .b(in[118]),
 .c(tree_684)
);
wire [0:0] tree_685;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_877 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[25]),
 .b(in[104]),
 .c(tree_685)
);
wire [0:0] tree_686;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_878 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[41]),
 .b(in[162]),
 .c(tree_686)
);
wire [0:0] tree_687;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_879 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[99]),
 .b(in[178]),
 .c(tree_687)
);
wire [0:0] tree_688;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_880 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_266),
 .b(tree_123),
 .c(tree_688)
);
wire [0:0] tree_689;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_881 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[52]),
 .b(in[129]),
 .c(tree_689)
);
wire [0:0] tree_690;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_882 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[101]),
 .b(in[147]),
 .c(tree_690)
);
wire [0:0] tree_691;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_883 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[73]),
 .b(1'h0),
 .c(tree_691)
);
wire [0:0] tree_692;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_884 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_691),
 .b(tree_6),
 .c(tree_692)
);
wire [0:0] tree_693;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_885 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[101]),
 .b(1'h0),
 .c(tree_693)
);
wire [0:0] tree_694;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_886 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_693),
 .b(tree_7),
 .c(tree_694)
);
wire [0:0] tree_695;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_887 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[85]),
 .b(1'h0),
 .c(tree_695)
);
wire [0:0] tree_696;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_888 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_695),
 .b(tree_9),
 .c(tree_696)
);
wire [0:0] tree_697;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_889 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[69]),
 .b(1'h0),
 .c(tree_697)
);
wire [0:0] tree_698;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_890 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_697),
 .b(tree_10),
 .c(tree_698)
);
wire [0:0] tree_699;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_891 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[160]),
 .b(1'h0),
 .c(tree_699)
);
wire [0:0] tree_700;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_892 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_699),
 .b(tree_14),
 .c(tree_700)
);
wire [0:0] tree_701;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_893 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_15),
 .b(tree_16),
 .c(tree_701)
);
wire [0:0] tree_702;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_894 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[176]),
 .b(1'h0),
 .c(tree_702)
);
wire [0:0] tree_703;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_895 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_702),
 .b(tree_21),
 .c(tree_703)
);
wire [0:0] tree_704;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_896 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_23),
 .b(tree_24),
 .c(tree_704)
);
wire [0:0] tree_705;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_897 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[152]),
 .b(1'h0),
 .c(tree_705)
);
wire [0:0] tree_706;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_898 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_705),
 .b(tree_26),
 .c(tree_706)
);
wire [0:0] tree_707;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_899 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_28),
 .b(tree_29),
 .c(tree_707)
);
wire [0:0] tree_708;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_900 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[8]),
 .b(1'h0),
 .c(tree_708)
);
wire [0:0] tree_709;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_901 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_708),
 .b(tree_30),
 .c(tree_709)
);
wire [0:0] tree_710;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_902 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[191]),
 .b(1'h0),
 .c(tree_710)
);
wire [0:0] tree_711;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_903 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_710),
 .b(tree_35),
 .c(tree_711)
);
wire [0:0] tree_712;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_904 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[126]),
 .b(1'h0),
 .c(tree_712)
);
wire [0:0] tree_713;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_905 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_712),
 .b(tree_38),
 .c(tree_713)
);
wire [0:0] tree_714;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_906 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[144]),
 .b(1'h0),
 .c(tree_714)
);
wire [0:0] tree_715;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_907 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_714),
 .b(tree_39),
 .c(tree_715)
);
wire [0:0] tree_716;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_908 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_40),
 .b(tree_41),
 .c(tree_716)
);
wire [0:0] tree_717;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_909 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[1]),
 .b(1'h0),
 .c(tree_717)
);
wire [0:0] tree_718;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_910 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_717),
 .b(tree_42),
 .c(tree_718)
);
wire [0:0] tree_719;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_911 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[13]),
 .b(1'h0),
 .c(tree_719)
);
wire [0:0] tree_720;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_912 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_719),
 .b(tree_43),
 .c(tree_720)
);
wire [0:0] tree_721;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_913 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[75]),
 .b(1'h0),
 .c(tree_721)
);
wire [0:0] tree_722;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_914 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_721),
 .b(tree_44),
 .c(tree_722)
);
wire [0:0] tree_723;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_915 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[118]),
 .b(1'h0),
 .c(tree_723)
);
wire [0:0] tree_724;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_916 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_723),
 .b(tree_46),
 .c(tree_724)
);
wire [0:0] tree_725;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_917 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[187]),
 .b(1'h0),
 .c(tree_725)
);
wire [0:0] tree_726;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_918 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_725),
 .b(tree_47),
 .c(tree_726)
);
wire [0:0] tree_727;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_919 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_48),
 .b(tree_49),
 .c(tree_727)
);
wire [0:0] tree_728;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_920 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[143]),
 .b(1'h0),
 .c(tree_728)
);
wire [0:0] tree_729;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_921 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_728),
 .b(tree_51),
 .c(tree_729)
);
wire [0:0] tree_730;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_922 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[170]),
 .b(1'h0),
 .c(tree_730)
);
wire [0:0] tree_731;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_923 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_730),
 .b(tree_53),
 .c(tree_731)
);
wire [0:0] tree_732;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_924 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[158]),
 .b(1'h0),
 .c(tree_732)
);
wire [0:0] tree_733;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_925 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_732),
 .b(tree_55),
 .c(tree_733)
);
wire [0:0] tree_734;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_926 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_56),
 .b(tree_57),
 .c(tree_734)
);
wire [0:0] tree_735;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_927 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2),
 .b(tree_59),
 .c(tree_735)
);
wire [0:0] tree_736;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_928 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_61),
 .b(tree_62),
 .c(tree_736)
);
wire [0:0] tree_737;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_929 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[133]),
 .b(1'h0),
 .c(tree_737)
);
wire [0:0] tree_738;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_930 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_737),
 .b(tree_64),
 .c(tree_738)
);
wire [0:0] tree_739;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_931 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_68),
 .b(tree_69),
 .c(tree_739)
);
wire [0:0] tree_740;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_932 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_70),
 .b(tree_32),
 .c(tree_740)
);
wire [0:0] tree_741;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_933 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_71),
 .b(tree_72),
 .c(tree_741)
);
wire [0:0] tree_742;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_934 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[74]),
 .b(1'h0),
 .c(tree_742)
);
wire [0:0] tree_743;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_935 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_742),
 .b(tree_73),
 .c(tree_743)
);
wire [0:0] tree_744;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_936 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[124]),
 .b(1'h0),
 .c(tree_744)
);
wire [0:0] tree_745;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_937 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_744),
 .b(tree_74),
 .c(tree_745)
);
wire [0:0] tree_746;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_938 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[150]),
 .b(1'h0),
 .c(tree_746)
);
wire [0:0] tree_747;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_939 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_746),
 .b(tree_76),
 .c(tree_747)
);
wire [0:0] tree_748;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_940 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[154]),
 .b(1'h0),
 .c(tree_748)
);
wire [0:0] tree_749;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_941 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_748),
 .b(tree_77),
 .c(tree_749)
);
wire [0:0] tree_750;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_942 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[78]),
 .b(1'h0),
 .c(tree_750)
);
wire [0:0] tree_751;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_943 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_750),
 .b(tree_78),
 .c(tree_751)
);
wire [0:0] tree_752;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_944 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[185]),
 .b(1'h0),
 .c(tree_752)
);
wire [0:0] tree_753;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_945 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_752),
 .b(tree_81),
 .c(tree_753)
);
wire [0:0] tree_754;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_946 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[65]),
 .b(1'h0),
 .c(tree_754)
);
wire [0:0] tree_755;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_947 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_754),
 .b(tree_82),
 .c(tree_755)
);
wire [0:0] tree_756;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_948 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_84),
 .b(tree_85),
 .c(tree_756)
);
wire [0:0] tree_757;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_949 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[87]),
 .b(1'h0),
 .c(tree_757)
);
wire [0:0] tree_758;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_950 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_757),
 .b(tree_86),
 .c(tree_758)
);
wire [0:0] tree_759;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_951 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[114]),
 .b(1'h0),
 .c(tree_759)
);
wire [0:0] tree_760;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_952 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_759),
 .b(tree_87),
 .c(tree_760)
);
wire [0:0] tree_761;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_953 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_58),
 .b(1'h0),
 .c(tree_761)
);
wire [0:0] tree_762;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_954 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_761),
 .b(tree_735),
 .c(tree_762)
);
wire [0:0] tree_763;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_955 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[63]),
 .b(1'h0),
 .c(tree_763)
);
wire [0:0] tree_764;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_956 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_763),
 .b(tree_88),
 .c(tree_764)
);
wire [0:0] tree_765;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_957 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[172]),
 .b(1'h0),
 .c(tree_765)
);
wire [0:0] tree_766;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_958 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_765),
 .b(tree_89),
 .c(tree_766)
);
wire [0:0] tree_767;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_959 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[128]),
 .b(1'h0),
 .c(tree_767)
);
wire [0:0] tree_768;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_960 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_767),
 .b(tree_91),
 .c(tree_768)
);
wire [0:0] tree_769;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_961 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[175]),
 .b(1'h0),
 .c(tree_769)
);
wire [0:0] tree_770;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_962 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_769),
 .b(1'h0),
 .c(tree_770)
);
wire [0:0] tree_771;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_963 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_770),
 .b(tree_95),
 .c(tree_771)
);
wire [0:0] tree_772;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_964 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[179]),
 .b(1'h0),
 .c(tree_772)
);
wire [0:0] tree_773;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_965 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_772),
 .b(tree_96),
 .c(tree_773)
);
wire [0:0] tree_774;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_966 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_38),
 .b(tree_97),
 .c(tree_774)
);
wire [0:0] tree_775;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_967 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_55),
 .b(tree_98),
 .c(tree_775)
);
wire [0:0] tree_776;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_968 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[188]),
 .b(1'h0),
 .c(tree_776)
);
wire [0:0] tree_777;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_969 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_776),
 .b(tree_99),
 .c(tree_777)
);
wire [0:0] tree_778;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_970 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[164]),
 .b(1'h0),
 .c(tree_778)
);
wire [0:0] tree_779;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_971 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_778),
 .b(tree_100),
 .c(tree_779)
);
wire [0:0] tree_780;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_972 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_101),
 .b(tree_102),
 .c(tree_780)
);
wire [0:0] tree_781;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_973 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[61]),
 .b(1'h0),
 .c(tree_781)
);
wire [0:0] tree_782;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_974 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_781),
 .b(tree_107),
 .c(tree_782)
);
wire [0:0] tree_783;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_975 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[43]),
 .b(1'h0),
 .c(tree_783)
);
wire [0:0] tree_784;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_976 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_783),
 .b(tree_108),
 .c(tree_784)
);
wire [0:0] tree_785;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_977 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[174]),
 .b(1'h0),
 .c(tree_785)
);
wire [0:0] tree_786;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_978 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_785),
 .b(tree_111),
 .c(tree_786)
);
wire [0:0] tree_787;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_979 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[182]),
 .b(1'h0),
 .c(tree_787)
);
wire [0:0] tree_788;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_980 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_787),
 .b(1'h0),
 .c(tree_788)
);
wire [0:0] tree_789;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_981 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_788),
 .b(tree_116),
 .c(tree_789)
);
wire [0:0] tree_790;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_982 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_9),
 .b(tree_117),
 .c(tree_790)
);
wire [0:0] tree_791;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_983 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_118),
 .b(tree_119),
 .c(tree_791)
);
wire [0:0] tree_792;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_984 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_120),
 .b(tree_121),
 .c(tree_792)
);
wire [0:0] tree_793;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_985 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_68),
 .b(1'h0),
 .c(tree_793)
);
wire [0:0] tree_794;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_986 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_793),
 .b(tree_694),
 .c(tree_794)
);
wire [0:0] tree_795;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_987 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[104]),
 .b(1'h0),
 .c(tree_795)
);
wire [0:0] tree_796;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_988 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_795),
 .b(tree_126),
 .c(tree_796)
);
wire [0:0] tree_797;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_989 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[10]),
 .b(1'h0),
 .c(tree_797)
);
wire [0:0] tree_798;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_990 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_797),
 .b(tree_129),
 .c(tree_798)
);
wire [0:0] tree_799;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_991 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[156]),
 .b(1'h0),
 .c(tree_799)
);
wire [0:0] tree_800;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_992 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_799),
 .b(tree_132),
 .c(tree_800)
);
wire [0:0] tree_801;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_993 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[41]),
 .b(1'h0),
 .c(tree_801)
);
wire [0:0] tree_802;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_994 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_801),
 .b(tree_133),
 .c(tree_802)
);
wire [0:0] tree_803;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_995 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[110]),
 .b(1'h0),
 .c(tree_803)
);
wire [0:0] tree_804;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_996 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_803),
 .b(tree_136),
 .c(tree_804)
);
wire [0:0] tree_805;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_997 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[191]),
 .b(1'h0),
 .c(tree_805)
);
wire [0:0] tree_806;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_998 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_805),
 .b(tree_137),
 .c(tree_806)
);
wire [0:0] tree_807;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_999 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_138),
 .b(tree_18),
 .c(tree_807)
);
wire [0:0] tree_808;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1000 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_139),
 .b(tree_140),
 .c(tree_808)
);
wire [0:0] tree_809;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1001 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_141),
 .b(tree_118),
 .c(tree_809)
);
wire [0:0] tree_810;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1002 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_144),
 .b(tree_145),
 .c(tree_810)
);
wire [0:0] tree_811;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1003 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_4),
 .b(tree_147),
 .c(tree_811)
);
wire [0:0] tree_812;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1004 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_150),
 .b(1'h0),
 .c(tree_812)
);
wire [0:0] tree_813;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1005 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_812),
 .b(tree_149),
 .c(tree_813)
);
wire [0:0] tree_814;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1006 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_51),
 .b(tree_156),
 .c(tree_814)
);
wire [0:0] tree_815;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1007 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_157),
 .b(tree_158),
 .c(tree_815)
);
wire [0:0] tree_816;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1008 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[45]),
 .b(1'h0),
 .c(tree_816)
);
wire [0:0] tree_817;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1009 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_816),
 .b(tree_159),
 .c(tree_817)
);
wire [0:0] tree_818;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1010 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_160),
 .b(tree_139),
 .c(tree_818)
);
wire [0:0] tree_819;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1011 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[29]),
 .b(1'h0),
 .c(tree_819)
);
wire [0:0] tree_820;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1012 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_819),
 .b(1'h0),
 .c(tree_820)
);
wire [0:0] tree_821;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1013 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_820),
 .b(tree_751),
 .c(tree_821)
);
wire [0:0] tree_822;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1014 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[49]),
 .b(1'h0),
 .c(tree_822)
);
wire [0:0] tree_823;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1015 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_822),
 .b(tree_161),
 .c(tree_823)
);
wire [0:0] tree_824;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1016 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_96),
 .b(tree_162),
 .c(tree_824)
);
wire [0:0] tree_825;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1017 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_0),
 .b(tree_163),
 .c(tree_825)
);
wire [0:0] tree_826;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1018 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_164),
 .b(1'h0),
 .c(tree_826)
);
wire [0:0] tree_827;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1019 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_826),
 .b(tree_149),
 .c(tree_827)
);
wire [0:0] tree_828;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1020 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[139]),
 .b(1'h0),
 .c(tree_828)
);
wire [0:0] tree_829;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1021 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_828),
 .b(tree_165),
 .c(tree_829)
);
wire [0:0] tree_830;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1022 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_166),
 .b(tree_167),
 .c(tree_830)
);
wire [0:0] tree_831;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1023 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[16]),
 .b(1'h0),
 .c(tree_831)
);
wire [0:0] tree_832;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1024 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_831),
 .b(tree_168),
 .c(tree_832)
);
wire [0:0] tree_833;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1025 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_170),
 .b(1'h0),
 .c(tree_833)
);
wire [0:0] tree_834;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1026 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_833),
 .b(tree_753),
 .c(tree_834)
);
wire [0:0] tree_835;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1027 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[146]),
 .b(1'h0),
 .c(tree_835)
);
wire [0:0] tree_836;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1028 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_835),
 .b(tree_173),
 .c(tree_836)
);
wire [0:0] tree_837;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1029 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[81]),
 .b(1'h0),
 .c(tree_837)
);
wire [0:0] tree_838;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1030 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_837),
 .b(1'h0),
 .c(tree_838)
);
wire [0:0] tree_839;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1031 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_838),
 .b(tree_177),
 .c(tree_839)
);
wire [0:0] tree_840;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1032 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_78),
 .b(1'h0),
 .c(tree_840)
);
wire [0:0] tree_841;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1033 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_840),
 .b(tree_729),
 .c(tree_841)
);
wire [0:0] tree_842;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1034 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_180),
 .b(tree_62),
 .c(tree_842)
);
wire [0:0] tree_843;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1035 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[70]),
 .b(1'h0),
 .c(tree_843)
);
wire [0:0] tree_844;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1036 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_843),
 .b(tree_182),
 .c(tree_844)
);
wire [0:0] tree_845;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1037 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_28),
 .b(tree_184),
 .c(tree_845)
);
wire [0:0] tree_846;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1038 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_185),
 .b(1'h0),
 .c(tree_846)
);
wire [0:0] tree_847;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1039 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_846),
 .b(tree_187),
 .c(tree_847)
);
wire [0:0] tree_848;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1040 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_189),
 .b(tree_163),
 .c(tree_848)
);
wire [0:0] tree_849;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1041 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[74]),
 .b(1'h0),
 .c(tree_849)
);
wire [0:0] tree_850;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1042 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_849),
 .b(tree_193),
 .c(tree_850)
);
wire [0:0] tree_851;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1043 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[138]),
 .b(1'h0),
 .c(tree_851)
);
wire [0:0] tree_852;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1044 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_851),
 .b(tree_194),
 .c(tree_852)
);
wire [0:0] tree_853;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1045 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_189),
 .b(tree_195),
 .c(tree_853)
);
wire [0:0] tree_854;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1046 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[102]),
 .b(1'h0),
 .c(tree_854)
);
wire [0:0] tree_855;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1047 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_854),
 .b(tree_198),
 .c(tree_855)
);
wire [0:0] tree_856;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1048 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_78),
 .b(tree_201),
 .c(tree_856)
);
wire [0:0] tree_857;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1049 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_84),
 .b(tree_202),
 .c(tree_857)
);
wire [0:0] tree_858;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1050 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_205),
 .b(tree_206),
 .c(tree_858)
);
wire [0:0] tree_859;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1051 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_101),
 .b(1'h0),
 .c(tree_859)
);
wire [0:0] tree_860;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1052 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_859),
 .b(tree_208),
 .c(tree_860)
);
wire [0:0] tree_861;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1053 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_209),
 .b(tree_210),
 .c(tree_861)
);
wire [0:0] tree_862;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1054 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[184]),
 .b(1'h0),
 .c(tree_862)
);
wire [0:0] tree_863;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1055 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_862),
 .b(tree_212),
 .c(tree_863)
);
wire [0:0] tree_864;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1056 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[173]),
 .b(1'h0),
 .c(tree_864)
);
wire [0:0] tree_865;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1057 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_864),
 .b(tree_221),
 .c(tree_865)
);
wire [0:0] tree_866;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1058 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[30]),
 .b(1'h0),
 .c(tree_866)
);
wire [0:0] tree_867;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1059 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_866),
 .b(tree_222),
 .c(tree_867)
);
wire [0:0] tree_868;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1060 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[131]),
 .b(1'h0),
 .c(tree_868)
);
wire [0:0] tree_869;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1061 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_868),
 .b(1'h0),
 .c(tree_869)
);
wire [0:0] tree_870;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1062 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_869),
 .b(tree_224),
 .c(tree_870)
);
wire [0:0] tree_871;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1063 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[187]),
 .b(1'h0),
 .c(tree_871)
);
wire [0:0] tree_872;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1064 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_871),
 .b(tree_225),
 .c(tree_872)
);
wire [0:0] tree_873;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1065 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_226),
 .b(tree_227),
 .c(tree_873)
);
wire [0:0] tree_874;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1066 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_98),
 .b(tree_228),
 .c(tree_874)
);
wire [0:0] tree_875;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1067 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_231),
 .b(1'h0),
 .c(tree_875)
);
wire [0:0] tree_876;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1068 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_875),
 .b(tree_230),
 .c(tree_876)
);
wire [0:0] tree_877;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1069 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_105),
 .b(1'h0),
 .c(tree_877)
);
wire [0:0] tree_878;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1070 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_877),
 .b(tree_707),
 .c(tree_878)
);
wire [0:0] tree_879;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1071 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[171]),
 .b(1'h0),
 .c(tree_879)
);
wire [0:0] tree_880;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1072 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_879),
 .b(1'h0),
 .c(tree_880)
);
wire [0:0] tree_881;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1073 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_880),
 .b(tree_238),
 .c(tree_881)
);
wire [0:0] tree_882;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1074 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_245),
 .b(tree_34),
 .c(tree_882)
);
wire [0:0] tree_883;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1075 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_171),
 .b(1'h0),
 .c(tree_883)
);
wire [0:0] tree_884;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1076 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_883),
 .b(tree_800),
 .c(tree_884)
);
wire [0:0] tree_885;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1077 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_123),
 .b(1'h0),
 .c(tree_885)
);
wire [0:0] tree_886;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1078 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_885),
 .b(tree_692),
 .c(tree_886)
);
wire [0:0] tree_887;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1079 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_247),
 .b(tree_248),
 .c(tree_887)
);
wire [0:0] tree_888;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1080 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_249),
 .b(tree_250),
 .c(tree_888)
);
wire [0:0] tree_889;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1081 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_46),
 .b(tree_252),
 .c(tree_889)
);
wire [0:0] tree_890;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1082 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[65]),
 .b(1'h0),
 .c(tree_890)
);
wire [0:0] tree_891;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1083 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_890),
 .b(tree_260),
 .c(tree_891)
);
wire [0:0] tree_892;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1084 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_263),
 .b(tree_264),
 .c(tree_892)
);
wire [0:0] tree_893;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1085 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_249),
 .b(tree_265),
 .c(tree_893)
);
wire [0:0] tree_894;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1086 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[121]),
 .b(1'h0),
 .c(tree_894)
);
wire [0:0] tree_895;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1087 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_894),
 .b(tree_266),
 .c(tree_895)
);
wire [0:0] tree_896;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1088 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[177]),
 .b(1'h0),
 .c(tree_896)
);
wire [0:0] tree_897;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1089 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_896),
 .b(tree_270),
 .c(tree_897)
);
wire [0:0] tree_898;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1090 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[169]),
 .b(1'h0),
 .c(tree_898)
);
wire [0:0] tree_899;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1091 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_898),
 .b(tree_274),
 .c(tree_899)
);
wire [0:0] tree_900;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1092 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[13]),
 .b(1'h0),
 .c(tree_900)
);
wire [0:0] tree_901;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1093 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_900),
 .b(1'h0),
 .c(tree_901)
);
wire [0:0] tree_902;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1094 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_901),
 .b(tree_782),
 .c(tree_902)
);
wire [0:0] tree_903;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1095 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[87]),
 .b(1'h0),
 .c(tree_903)
);
wire [0:0] tree_904;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1096 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_903),
 .b(1'h0),
 .c(tree_904)
);
wire [0:0] tree_905;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1097 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_904),
 .b(tree_798),
 .c(tree_905)
);
wire [0:0] tree_906;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1098 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[184]),
 .b(1'h0),
 .c(tree_906)
);
wire [0:0] tree_907;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1099 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_906),
 .b(tree_275),
 .c(tree_907)
);
wire [0:0] tree_908;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1100 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_277),
 .b(tree_278),
 .c(tree_908)
);
wire [0:0] tree_909;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1101 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_279),
 .b(tree_280),
 .c(tree_909)
);
wire [0:0] tree_910;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1102 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_281),
 .b(1'h0),
 .c(tree_910)
);
wire [0:0] tree_911;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1103 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_910),
 .b(tree_701),
 .c(tree_911)
);
wire [0:0] tree_912;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1104 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_73),
 .b(1'h0),
 .c(tree_912)
);
wire [0:0] tree_913;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1105 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_912),
 .b(tree_284),
 .c(tree_913)
);
wire [0:0] tree_914;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1106 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[120]),
 .b(1'h0),
 .c(tree_914)
);
wire [0:0] tree_915;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1107 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_914),
 .b(tree_285),
 .c(tree_915)
);
wire [0:0] tree_916;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1108 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[44]),
 .b(1'h0),
 .c(tree_916)
);
wire [0:0] tree_917;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1109 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_916),
 .b(tree_299),
 .c(tree_917)
);
wire [0:0] tree_918;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1110 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[50]),
 .b(1'h0),
 .c(tree_918)
);
wire [0:0] tree_919;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1111 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_918),
 .b(1'h0),
 .c(tree_919)
);
wire [0:0] tree_920;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1112 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_919),
 .b(tree_711),
 .c(tree_920)
);
wire [0:0] tree_921;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1113 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_5),
 .b(tree_302),
 .c(tree_921)
);
wire [0:0] tree_922;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1114 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_304),
 .b(tree_709),
 .c(tree_922)
);
wire [0:0] tree_923;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1115 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[29]),
 .b(1'h0),
 .c(tree_923)
);
wire [0:0] tree_924;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1116 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_923),
 .b(tree_305),
 .c(tree_924)
);
wire [0:0] tree_925;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1117 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_307),
 .b(tree_309),
 .c(tree_925)
);
wire [0:0] tree_926;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1118 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[36]),
 .b(1'h0),
 .c(tree_926)
);
wire [0:0] tree_927;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1119 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_926),
 .b(tree_311),
 .c(tree_927)
);
wire [0:0] tree_928;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1120 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[72]),
 .b(1'h0),
 .c(tree_928)
);
wire [0:0] tree_929;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1121 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_928),
 .b(tree_319),
 .c(tree_929)
);
wire [0:0] tree_930;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1122 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_167),
 .b(tree_321),
 .c(tree_930)
);
wire [0:0] tree_931;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1123 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_271),
 .b(tree_322),
 .c(tree_931)
);
wire [0:0] tree_932;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1124 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_252),
 .b(tree_327),
 .c(tree_932)
);
wire [0:0] tree_933;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1125 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_138),
 .b(1'h0),
 .c(tree_933)
);
wire [0:0] tree_934;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1126 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_933),
 .b(tree_696),
 .c(tree_934)
);
wire [0:0] tree_935;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1127 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_209),
 .b(tree_330),
 .c(tree_935)
);
wire [0:0] tree_936;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1128 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[113]),
 .b(1'h0),
 .c(tree_936)
);
wire [0:0] tree_937;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1129 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_936),
 .b(tree_331),
 .c(tree_937)
);
wire [0:0] tree_938;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1130 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_836),
 .b(tree_110),
 .c(tree_938)
);
wire [0:0] tree_939;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1131 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[143]),
 .b(1'h0),
 .c(tree_939)
);
wire [0:0] tree_940;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1132 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_939),
 .b(tree_334),
 .c(tree_940)
);
wire [0:0] tree_941;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1133 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[129]),
 .b(1'h0),
 .c(tree_941)
);
wire [0:0] tree_942;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1134 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_941),
 .b(tree_335),
 .c(tree_942)
);
wire [0:0] tree_943;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1135 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[65]),
 .b(1'h0),
 .c(tree_943)
);
wire [0:0] tree_944;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1136 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_943),
 .b(tree_337),
 .c(tree_944)
);
wire [0:0] tree_945;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1137 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[169]),
 .b(1'h0),
 .c(tree_945)
);
wire [0:0] tree_946;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1138 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_945),
 .b(tree_339),
 .c(tree_946)
);
wire [0:0] tree_947;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1139 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_157),
 .b(tree_342),
 .c(tree_947)
);
wire [0:0] tree_948;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1140 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_344),
 .b(tree_346),
 .c(tree_948)
);
wire [0:0] tree_949;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1141 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_351),
 .b(tree_353),
 .c(tree_949)
);
wire [0:0] tree_950;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1142 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[115]),
 .b(1'h0),
 .c(tree_950)
);
wire [0:0] tree_951;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1143 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_950),
 .b(tree_358),
 .c(tree_951)
);
wire [0:0] tree_952;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1144 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[187]),
 .b(1'h0),
 .c(tree_952)
);
wire [0:0] tree_953;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1145 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_952),
 .b(tree_360),
 .c(tree_953)
);
wire [0:0] tree_954;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1146 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_361),
 .b(tree_362),
 .c(tree_954)
);
wire [0:0] tree_955;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1147 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[116]),
 .b(1'h0),
 .c(tree_955)
);
wire [0:0] tree_956;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1148 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_955),
 .b(1'h0),
 .c(tree_956)
);
wire [0:0] tree_957;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1149 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_956),
 .b(tree_364),
 .c(tree_957)
);
wire [0:0] tree_958;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1150 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_366),
 .b(1'h0),
 .c(tree_958)
);
wire [0:0] tree_959;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1151 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_958),
 .b(tree_815),
 .c(tree_959)
);
wire [0:0] tree_960;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1152 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[66]),
 .b(1'h0),
 .c(tree_960)
);
wire [0:0] tree_961;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1153 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_960),
 .b(tree_376),
 .c(tree_961)
);
wire [0:0] tree_962;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1154 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_378),
 .b(tree_379),
 .c(tree_962)
);
wire [0:0] tree_963;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1155 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_380),
 .b(1'h0),
 .c(tree_963)
);
wire [0:0] tree_964;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1156 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_963),
 .b(tree_382),
 .c(tree_964)
);
wire [0:0] tree_965;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1157 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[172]),
 .b(1'h0),
 .c(tree_965)
);
wire [0:0] tree_966;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1158 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_965),
 .b(tree_386),
 .c(tree_966)
);
wire [0:0] tree_967;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1159 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[189]),
 .b(1'h0),
 .c(tree_967)
);
wire [0:0] tree_968;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1160 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_967),
 .b(tree_392),
 .c(tree_968)
);
wire [0:0] tree_969;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1161 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_100),
 .b(tree_395),
 .c(tree_969)
);
wire [0:0] tree_970;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1162 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_354),
 .b(tree_396),
 .c(tree_970)
);
wire [0:0] tree_971;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1163 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_397),
 .b(1'h0),
 .c(tree_971)
);
wire [0:0] tree_972;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1164 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_971),
 .b(tree_304),
 .c(tree_972)
);
wire [0:0] tree_973;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1165 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_248),
 .b(1'h0),
 .c(tree_973)
);
wire [0:0] tree_974;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1166 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_973),
 .b(tree_399),
 .c(tree_974)
);
wire [0:0] tree_975;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1167 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_245),
 .b(tree_400),
 .c(tree_975)
);
wire [0:0] tree_976;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1168 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_412),
 .b(1'h0),
 .c(tree_976)
);
wire [0:0] tree_977;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1169 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_976),
 .b(tree_413),
 .c(tree_977)
);
wire [0:0] tree_978;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1170 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_426),
 .b(1'h0),
 .c(tree_978)
);
wire [0:0] tree_979;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1171 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_425),
 .b(tree_978),
 .c(tree_979)
);
wire [0:0] tree_980;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1172 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_428),
 .b(tree_429),
 .c(tree_980)
);
wire [0:0] tree_981;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1173 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[112]),
 .b(1'h0),
 .c(tree_981)
);
wire [0:0] tree_982;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1174 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_981),
 .b(1'h0),
 .c(tree_982)
);
wire [0:0] tree_983;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1175 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_982),
 .b(tree_430),
 .c(tree_983)
);
wire [0:0] tree_984;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1176 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[30]),
 .b(1'h0),
 .c(tree_984)
);
wire [0:0] tree_985;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1177 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_984),
 .b(1'h0),
 .c(tree_985)
);
wire [0:0] tree_986;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1178 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_985),
 .b(tree_915),
 .c(tree_986)
);
wire [0:0] tree_987;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1179 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[45]),
 .b(1'h0),
 .c(tree_987)
);
wire [0:0] tree_988;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1180 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_987),
 .b(1'h0),
 .c(tree_988)
);
wire [0:0] tree_989;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1181 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_988),
 .b(tree_889),
 .c(tree_989)
);
wire [0:0] tree_990;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1182 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_39),
 .b(tree_448),
 .c(tree_990)
);
wire [0:0] tree_991;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1183 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_460),
 .b(tree_461),
 .c(tree_991)
);
wire [0:0] tree_992;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1184 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[149]),
 .b(1'h0),
 .c(tree_992)
);
wire [0:0] tree_993;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1185 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_992),
 .b(tree_462),
 .c(tree_993)
);
wire [0:0] tree_994;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1186 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_111),
 .b(tree_463),
 .c(tree_994)
);
wire [0:0] tree_995;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1187 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_465),
 .b(1'h0),
 .c(tree_995)
);
wire [0:0] tree_996;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1188 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_995),
 .b(tree_777),
 .c(tree_996)
);
wire [0:0] tree_997;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1189 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_467),
 .b(tree_469),
 .c(tree_997)
);
wire [0:0] tree_998;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1190 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_48),
 .b(tree_471),
 .c(tree_998)
);
wire [0:0] tree_999;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1191 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[140]),
 .b(1'h0),
 .c(tree_999)
);
wire [0:0] tree_1000;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1192 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_999),
 .b(1'h0),
 .c(tree_1000)
);
wire [0:0] tree_1001;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1193 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1000),
 .b(tree_756),
 .c(tree_1001)
);
wire [0:0] tree_1002;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1194 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_453),
 .b(1'h0),
 .c(tree_1002)
);
wire [0:0] tree_1003;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1195 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_755),
 .b(tree_1002),
 .c(tree_1003)
);
wire [0:0] tree_1004;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1196 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_483),
 .b(1'h0),
 .c(tree_1004)
);
wire [0:0] tree_1005;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1197 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1004),
 .b(tree_230),
 .c(tree_1005)
);
wire [0:0] tree_1006;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1198 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[57]),
 .b(1'h0),
 .c(tree_1006)
);
wire [0:0] tree_1007;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1199 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1006),
 .b(1'h0),
 .c(tree_1007)
);
wire [0:0] tree_1008;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1200 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1007),
 .b(tree_694),
 .c(tree_1008)
);
wire [0:0] tree_1009;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1201 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_190),
 .b(tree_489),
 .c(tree_1009)
);
wire [0:0] tree_1010;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1202 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_490),
 .b(1'h0),
 .c(tree_1010)
);
wire [0:0] tree_1011;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1203 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_415),
 .b(tree_1010),
 .c(tree_1011)
);
wire [0:0] tree_1012;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1204 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[139]),
 .b(1'h0),
 .c(tree_1012)
);
wire [0:0] tree_1013;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1205 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1012),
 .b(1'h0),
 .c(tree_1013)
);
wire [0:0] tree_1014;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1206 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1013),
 .b(tree_494),
 .c(tree_1014)
);
wire [0:0] tree_1015;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1207 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_104),
 .b(tree_502),
 .c(tree_1015)
);
wire [0:0] tree_1016;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1208 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_402),
 .b(1'h0),
 .c(tree_1016)
);
wire [0:0] tree_1017;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1209 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1016),
 .b(tree_504),
 .c(tree_1017)
);
wire [0:0] tree_1018;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1210 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_506),
 .b(tree_507),
 .c(tree_1018)
);
wire [0:0] tree_1019;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1211 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_171),
 .b(1'h0),
 .c(tree_1019)
);
wire [0:0] tree_1020;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1212 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1019),
 .b(tree_515),
 .c(tree_1020)
);
wire [0:0] tree_1021;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1213 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[149]),
 .b(1'h0),
 .c(tree_1021)
);
wire [0:0] tree_1022;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1214 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1021),
 .b(1'h0),
 .c(tree_1022)
);
wire [0:0] tree_1023;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1215 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1022),
 .b(tree_975),
 .c(tree_1023)
);
wire [0:0] tree_1024;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1216 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_97),
 .b(1'h0),
 .c(tree_1024)
);
wire [0:0] tree_1025;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1217 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1024),
 .b(tree_525),
 .c(tree_1025)
);
wire [0:0] tree_1026;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1218 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_334),
 .b(1'h0),
 .c(tree_1026)
);
wire [0:0] tree_1027;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1219 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1026),
 .b(tree_541),
 .c(tree_1027)
);
wire [0:0] tree_1028;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1220 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_299),
 .b(tree_542),
 .c(tree_1028)
);
wire [0:0] tree_1029;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1221 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_40),
 .b(1'h0),
 .c(tree_1029)
);
wire [0:0] tree_1030;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1222 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1029),
 .b(tree_558),
 .c(tree_1030)
);
wire [0:0] tree_1031;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1223 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_397),
 .b(tree_559),
 .c(tree_1031)
);
wire [0:0] tree_1032;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1224 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_416),
 .b(1'h0),
 .c(tree_1032)
);
wire [0:0] tree_1033;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1225 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1032),
 .b(1'h0),
 .c(tree_1033)
);
wire [0:0] tree_1034;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1226 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1033),
 .b(tree_881),
 .c(tree_1034)
);
wire [0:0] tree_1035;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1227 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[114]),
 .b(1'h0),
 .c(tree_1035)
);
wire [0:0] tree_1036;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1228 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1035),
 .b(tree_583),
 .c(tree_1036)
);
wire [0:0] tree_1037;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1229 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_585),
 .b(tree_587),
 .c(tree_1037)
);
wire [0:0] tree_1038;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1230 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[125]),
 .b(1'h0),
 .c(tree_1038)
);
wire [0:0] tree_1039;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1231 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1038),
 .b(1'h0),
 .c(tree_1039)
);
wire [0:0] tree_1040;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1232 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1039),
 .b(tree_897),
 .c(tree_1040)
);
wire [0:0] tree_1041;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1233 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_542),
 .b(tree_596),
 .c(tree_1041)
);
wire [0:0] tree_1042;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1234 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_319),
 .b(tree_601),
 .c(tree_1042)
);
wire [0:0] tree_1043;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1235 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[84]),
 .b(in[12]),
 .c(tree_1043)
);
wire [0:0] tree_1044;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1236 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1043),
 .b(tree_85),
 .c(tree_1044)
);
wire [0:0] tree_1045;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1237 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_360),
 .b(tree_29),
 .c(tree_1045)
);
wire [0:0] tree_1046;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1238 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_39),
 .b(tree_158),
 .c(tree_1046)
);
wire [0:0] tree_1047;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1239 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_572),
 .b(tree_559),
 .c(tree_1047)
);
wire [0:0] tree_1048;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1240 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_606),
 .b(tree_603),
 .c(tree_1048)
);
wire [0:0] tree_1049;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1241 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1044),
 .b(tree_1045),
 .c(tree_1049)
);
wire [0:0] tree_1050;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1242 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1046),
 .b(tree_1047),
 .c(tree_1050)
);
wire [0:0] tree_1051;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1243 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1048),
 .b(tree_915),
 .c(tree_1051)
);
wire [0:0] tree_1052;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1244 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_95),
 .b(tree_494),
 .c(tree_1052)
);
wire [0:0] tree_1053;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1245 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_598),
 .b(tree_718),
 .c(tree_1053)
);
wire [0:0] tree_1054;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1246 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_722),
 .b(tree_605),
 .c(tree_1054)
);
wire [0:0] tree_1055;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1247 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_608),
 .b(tree_574),
 .c(tree_1055)
);
wire [0:0] tree_1056;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1248 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_488),
 .b(tree_423),
 .c(tree_1056)
);
wire [0:0] tree_1057;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1249 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_609),
 .b(tree_792),
 .c(tree_1057)
);
wire [0:0] tree_1058;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1250 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_610),
 .b(tree_432),
 .c(tree_1058)
);
wire [0:0] tree_1059;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1251 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1049),
 .b(tree_1050),
 .c(tree_1059)
);
wire [0:0] tree_1060;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1252 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1051),
 .b(tree_1052),
 .c(tree_1060)
);
wire [0:0] tree_1061;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1253 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1053),
 .b(tree_1054),
 .c(tree_1061)
);
wire [0:0] tree_1062;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1254 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1055),
 .b(tree_1056),
 .c(tree_1062)
);
wire [0:0] tree_1063;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1255 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1057),
 .b(tree_1058),
 .c(tree_1063)
);
wire [0:0] tree_1064;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1256 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_529),
 .b(tree_1023),
 .c(tree_1064)
);
wire [0:0] tree_1065;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1257 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_870),
 .b(1'h0),
 .c(tree_1065)
);
wire [0:0] tree_1066;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1258 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1059),
 .b(tree_1060),
 .c(tree_1066)
);
wire [0:0] tree_1067;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1259 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1061),
 .b(tree_1062),
 .c(tree_1067)
);
wire [0:0] tree_1068;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1260 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1063),
 .b(tree_1064),
 .c(tree_1068)
);
wire [0:0] tree_1069;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1261 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1065),
 .b(1'h0),
 .c(tree_1069)
);
wire [0:0] tree_1070;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1262 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1066),
 .b(tree_1067),
 .c(tree_1070)
);
wire [0:0] tree_1071;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1263 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1068),
 .b(tree_1069),
 .c(tree_1071)
);
wire [0:0] tree_1072;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1264 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1070),
 .b(tree_1071),
 .c(tree_1072)
);
wire [0:0] tree_1073;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1265 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[49]),
 .b(in[121]),
 .c(tree_1073)
);
wire [0:0] tree_1074;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1266 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[147]),
 .b(in[149]),
 .c(tree_1074)
);
wire [0:0] tree_1075;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1267 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[150]),
 .b(1'h0),
 .c(tree_1075)
);
wire [0:0] tree_1076;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1268 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1073),
 .b(tree_1074),
 .c(tree_1076)
);
wire [0:0] tree_1077;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1269 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_39),
 .b(tree_1075),
 .c(tree_1077)
);
wire [0:0] tree_1078;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1270 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_62),
 .b(tree_55),
 .c(tree_1078)
);
wire [0:0] tree_1079;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1271 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_209),
 .b(tree_195),
 .c(tree_1079)
);
wire [0:0] tree_1080;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1272 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_80),
 .b(tree_323),
 .c(tree_1080)
);
wire [0:0] tree_1081;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1273 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_614),
 .b(tree_280),
 .c(tree_1081)
);
wire [0:0] tree_1082;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1274 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_20),
 .b(1'h0),
 .c(tree_1082)
);
wire [0:0] tree_1083;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1275 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1076),
 .b(tree_1077),
 .c(tree_1083)
);
wire [0:0] tree_1084;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1276 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1079),
 .b(tree_1078),
 .c(tree_1084)
);
wire [0:0] tree_1085;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1277 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1081),
 .b(tree_1080),
 .c(tree_1085)
);
wire [0:0] tree_1086;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1278 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1082),
 .b(tree_764),
 .c(tree_1086)
);
wire [0:0] tree_1087;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1279 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_546),
 .b(tree_612),
 .c(tree_1087)
);
wire [0:0] tree_1088;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1280 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_473),
 .b(tree_442),
 .c(tree_1088)
);
wire [0:0] tree_1089;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1281 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_932),
 .b(tree_307),
 .c(tree_1089)
);
wire [0:0] tree_1090;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1282 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_613),
 .b(tree_616),
 .c(tree_1090)
);
wire [0:0] tree_1091;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1283 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_824),
 .b(tree_618),
 .c(tree_1091)
);
wire [0:0] tree_1092;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1284 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1083),
 .b(tree_1084),
 .c(tree_1092)
);
wire [0:0] tree_1093;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1285 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1085),
 .b(tree_1086),
 .c(tree_1093)
);
wire [0:0] tree_1094;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1286 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1087),
 .b(tree_1088),
 .c(tree_1094)
);
wire [0:0] tree_1095;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1287 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1089),
 .b(tree_1090),
 .c(tree_1095)
);
wire [0:0] tree_1096;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1288 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1091),
 .b(tree_886),
 .c(tree_1096)
);
wire [0:0] tree_1097;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1289 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_876),
 .b(1'h0),
 .c(tree_1097)
);
wire [0:0] tree_1098;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1290 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1092),
 .b(tree_1093),
 .c(tree_1098)
);
wire [0:0] tree_1099;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1291 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1094),
 .b(tree_1095),
 .c(tree_1099)
);
wire [0:0] tree_1100;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1292 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1096),
 .b(tree_1097),
 .c(tree_1100)
);
wire [0:0] tree_1101;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1293 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1098),
 .b(tree_1099),
 .c(tree_1101)
);
wire [0:0] tree_1102;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1294 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1100),
 .b(1'h0),
 .c(tree_1102)
);
wire [0:0] tree_1103;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1295 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1101),
 .b(tree_1102),
 .c(tree_1103)
);
wire [0:0] tree_1104;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1296 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_144),
 .b(tree_622),
 .c(tree_1104)
);
wire [0:0] tree_1105;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1297 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[55]),
 .b(1'h0),
 .c(tree_1105)
);
wire [0:0] tree_1106;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1298 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1105),
 .b(1'h0),
 .c(tree_1106)
);
wire [0:0] tree_1107;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1299 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1106),
 .b(1'h0),
 .c(tree_1107)
);
wire [0:0] tree_1108;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1300 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1107),
 .b(tree_1005),
 .c(tree_1108)
);
wire [0:0] tree_1109;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1301 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2),
 .b(1'h0),
 .c(tree_1109)
);
wire [0:0] tree_1110;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1302 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1109),
 .b(tree_848),
 .c(tree_1110)
);
wire [0:0] tree_1111;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1303 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_231),
 .b(1'h0),
 .c(tree_1111)
);
wire [0:0] tree_1112;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1304 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1111),
 .b(tree_628),
 .c(tree_1112)
);
wire [0:0] tree_1113;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1305 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_620),
 .b(tree_629),
 .c(tree_1113)
);
wire [0:0] tree_1114;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1306 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_603),
 .b(1'h0),
 .c(tree_1114)
);
wire [0:0] tree_1115;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1307 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1114),
 .b(tree_786),
 .c(tree_1115)
);
wire [0:0] tree_1116;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1308 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_572),
 .b(1'h0),
 .c(tree_1116)
);
wire [0:0] tree_1117;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1309 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1116),
 .b(tree_631),
 .c(tree_1117)
);
wire [0:0] tree_1118;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1310 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[142]),
 .b(in[96]),
 .c(tree_1118)
);
wire [0:0] tree_1119;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1311 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[156]),
 .b(1'h0),
 .c(tree_1119)
);
wire [0:0] tree_1120;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1312 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1118),
 .b(tree_1119),
 .c(tree_1120)
);
wire [0:0] tree_1121;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1313 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_165),
 .b(tree_96),
 .c(tree_1121)
);
wire [0:0] tree_1122;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1314 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_583),
 .b(tree_61),
 .c(tree_1122)
);
wire [0:0] tree_1123;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1315 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_260),
 .b(tree_544),
 .c(tree_1123)
);
wire [0:0] tree_1124;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1316 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_386),
 .b(tree_133),
 .c(tree_1124)
);
wire [0:0] tree_1125;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1317 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_593),
 .b(tree_237),
 .c(tree_1125)
);
wire [0:0] tree_1126;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1318 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_632),
 .b(tree_602),
 .c(tree_1126)
);
wire [0:0] tree_1127;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1319 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1120),
 .b(tree_1121),
 .c(tree_1127)
);
wire [0:0] tree_1128;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1320 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1122),
 .b(tree_1123),
 .c(tree_1128)
);
wire [0:0] tree_1129;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1321 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1124),
 .b(tree_1125),
 .c(tree_1129)
);
wire [0:0] tree_1130;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1322 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_975),
 .b(tree_1126),
 .c(tree_1130)
);
wire [0:0] tree_1131;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1323 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_546),
 .b(tree_863),
 .c(tree_1131)
);
wire [0:0] tree_1132;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1324 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_850),
 .b(tree_385),
 .c(tree_1132)
);
wire [0:0] tree_1133;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1325 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_296),
 .b(tree_511),
 .c(tree_1133)
);
wire [0:0] tree_1134;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1326 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_633),
 .b(1'h0),
 .c(tree_1134)
);
wire [0:0] tree_1135;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1327 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1127),
 .b(tree_1128),
 .c(tree_1135)
);
wire [0:0] tree_1136;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1328 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1129),
 .b(tree_1130),
 .c(tree_1136)
);
wire [0:0] tree_1137;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1329 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1131),
 .b(tree_1132),
 .c(tree_1137)
);
wire [0:0] tree_1138;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1330 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1133),
 .b(tree_1134),
 .c(tree_1138)
);
wire [0:0] tree_1139;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1331 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1110),
 .b(1'h0),
 .c(tree_1139)
);
wire [0:0] tree_1140;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1332 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1135),
 .b(tree_1136),
 .c(tree_1140)
);
wire [0:0] tree_1141;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1333 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1137),
 .b(tree_1138),
 .c(tree_1141)
);
wire [0:0] tree_1142;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1334 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1139),
 .b(1'h0),
 .c(tree_1142)
);
wire [0:0] tree_1143;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1335 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1140),
 .b(tree_1141),
 .c(tree_1143)
);
wire [0:0] tree_1144;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1336 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1142),
 .b(1'h0),
 .c(tree_1144)
);
wire [0:0] tree_1145;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1337 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1143),
 .b(tree_1144),
 .c(tree_1145)
);
wire [0:0] tree_1146;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1338 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[18]),
 .b(in[19]),
 .c(tree_1146)
);
wire [0:0] tree_1147;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1339 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[107]),
 .b(in[131]),
 .c(tree_1147)
);
wire [0:0] tree_1148;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1340 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1146),
 .b(tree_1147),
 .c(tree_1148)
);
wire [0:0] tree_1149;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1341 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_280),
 .b(tree_119),
 .c(tree_1149)
);
wire [0:0] tree_1150;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1342 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_150),
 .b(tree_410),
 .c(tree_1150)
);
wire [0:0] tree_1151;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1343 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_338),
 .b(tree_634),
 .c(tree_1151)
);
wire [0:0] tree_1152;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1344 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_320),
 .b(1'h0),
 .c(tree_1152)
);
wire [0:0] tree_1153;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1345 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1148),
 .b(tree_1149),
 .c(tree_1153)
);
wire [0:0] tree_1154;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1346 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1150),
 .b(tree_1151),
 .c(tree_1154)
);
wire [0:0] tree_1155;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1347 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_131),
 .b(tree_1152),
 .c(tree_1155)
);
wire [0:0] tree_1156;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1348 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_565),
 .b(tree_961),
 .c(tree_1156)
);
wire [0:0] tree_1157;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1349 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_636),
 .b(tree_487),
 .c(tree_1157)
);
wire [0:0] tree_1158;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1350 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_842),
 .b(tree_893),
 .c(tree_1158)
);
wire [0:0] tree_1159;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1351 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_638),
 .b(tree_609),
 .c(tree_1159)
);
wire [0:0] tree_1160;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1352 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_994),
 .b(tree_780),
 .c(tree_1160)
);
wire [0:0] tree_1161;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1353 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1153),
 .b(tree_1154),
 .c(tree_1161)
);
wire [0:0] tree_1162;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1354 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1155),
 .b(tree_1156),
 .c(tree_1162)
);
wire [0:0] tree_1163;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1355 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1157),
 .b(tree_1158),
 .c(tree_1163)
);
wire [0:0] tree_1164;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1356 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1159),
 .b(tree_1160),
 .c(tree_1164)
);
wire [0:0] tree_1165;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1357 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_626),
 .b(tree_878),
 .c(tree_1165)
);
wire [0:0] tree_1166;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1358 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_641),
 .b(tree_643),
 .c(tree_1166)
);
wire [0:0] tree_1167;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1359 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1161),
 .b(tree_1162),
 .c(tree_1167)
);
wire [0:0] tree_1168;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1360 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1163),
 .b(tree_1164),
 .c(tree_1168)
);
wire [0:0] tree_1169;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1361 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1165),
 .b(tree_1166),
 .c(tree_1169)
);
wire [0:0] tree_1170;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1362 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1167),
 .b(tree_1168),
 .c(tree_1170)
);
wire [0:0] tree_1171;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1363 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1169),
 .b(1'h0),
 .c(tree_1171)
);
wire [0:0] tree_1172;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1364 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1170),
 .b(tree_1171),
 .c(tree_1172)
);
wire [0:0] tree_1173;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1365 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[41]),
 .b(in[9]),
 .c(tree_1173)
);
wire [0:0] tree_1174;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1366 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[80]),
 .b(in[120]),
 .c(tree_1174)
);
wire [0:0] tree_1175;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1367 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1173),
 .b(tree_1174),
 .c(tree_1175)
);
wire [0:0] tree_1176;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1368 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_270),
 .b(tree_38),
 .c(tree_1176)
);
wire [0:0] tree_1177;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1369 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_164),
 .b(tree_44),
 .c(tree_1177)
);
wire [0:0] tree_1178;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1370 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_226),
 .b(tree_167),
 .c(tree_1178)
);
wire [0:0] tree_1179;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1371 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_279),
 .b(tree_67),
 .c(tree_1179)
);
wire [0:0] tree_1180;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1372 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1175),
 .b(tree_1176),
 .c(tree_1180)
);
wire [0:0] tree_1181;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1373 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1177),
 .b(tree_1178),
 .c(tree_1181)
);
wire [0:0] tree_1182;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1374 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1179),
 .b(tree_863),
 .c(tree_1182)
);
wire [0:0] tree_1183;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1375 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_645),
 .b(tree_698),
 .c(tree_1183)
);
wire [0:0] tree_1184;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1376 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_353),
 .b(tree_796),
 .c(tree_1184)
);
wire [0:0] tree_1185;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1377 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_501),
 .b(tree_966),
 .c(tree_1185)
);
wire [0:0] tree_1186;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1378 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_513),
 .b(tree_646),
 .c(tree_1186)
);
wire [0:0] tree_1187;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1379 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_522),
 .b(tree_648),
 .c(tree_1187)
);
wire [0:0] tree_1188;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1380 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_649),
 .b(1'h0),
 .c(tree_1188)
);
wire [0:0] tree_1189;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1381 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1180),
 .b(tree_1181),
 .c(tree_1189)
);
wire [0:0] tree_1190;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1382 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1182),
 .b(tree_1183),
 .c(tree_1190)
);
wire [0:0] tree_1191;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1383 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1185),
 .b(tree_1184),
 .c(tree_1191)
);
wire [0:0] tree_1192;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1384 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1186),
 .b(tree_1187),
 .c(tree_1192)
);
wire [0:0] tree_1193;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1385 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_957),
 .b(tree_1188),
 .c(tree_1193)
);
wire [0:0] tree_1194;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1386 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1189),
 .b(tree_1190),
 .c(tree_1194)
);
wire [0:0] tree_1195;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1387 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1191),
 .b(tree_1192),
 .c(tree_1195)
);
wire [0:0] tree_1196;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1388 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1193),
 .b(1'h0),
 .c(tree_1196)
);
wire [0:0] tree_1197;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1389 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1194),
 .b(tree_1195),
 .c(tree_1197)
);
wire [0:0] tree_1198;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1390 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1196),
 .b(1'h0),
 .c(tree_1198)
);
wire [0:0] tree_1199;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1391 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1197),
 .b(tree_1198),
 .c(tree_1199)
);
wire [0:0] tree_1200;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1392 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_334),
 .b(1'h0),
 .c(tree_1200)
);
wire [0:0] tree_1201;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1393 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1200),
 .b(tree_655),
 .c(tree_1201)
);
wire [0:0] tree_1202;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1394 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_760),
 .b(tree_560),
 .c(tree_1202)
);
wire [0:0] tree_1203;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1395 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_663),
 .b(tree_784),
 .c(tree_1203)
);
wire [0:0] tree_1204;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1396 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[17]),
 .b(in[48]),
 .c(tree_1204)
);
wire [0:0] tree_1205;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1397 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[93]),
 .b(in[137]),
 .c(tree_1205)
);
wire [0:0] tree_1206;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1398 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[142]),
 .b(in[154]),
 .c(tree_1206)
);
wire [0:0] tree_1207;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1399 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[164]),
 .b(in[157]),
 .c(tree_1207)
);
wire [0:0] tree_1208;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1400 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1204),
 .b(tree_1205),
 .c(tree_1208)
);
wire [0:0] tree_1209;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1401 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1206),
 .b(tree_1207),
 .c(tree_1209)
);
wire [0:0] tree_1210;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1402 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_88),
 .b(tree_80),
 .c(tree_1210)
);
wire [0:0] tree_1211;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1403 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_172),
 .b(tree_403),
 .c(tree_1211)
);
wire [0:0] tree_1212;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1404 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_606),
 .b(1'h0),
 .c(tree_1212)
);
wire [0:0] tree_1213;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1405 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1208),
 .b(tree_1209),
 .c(tree_1213)
);
wire [0:0] tree_1214;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1406 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1210),
 .b(tree_1211),
 .c(tree_1214)
);
wire [0:0] tree_1215;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1407 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1212),
 .b(tree_430),
 .c(tree_1215)
);
wire [0:0] tree_1216;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1408 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_287),
 .b(tree_628),
 .c(tree_1216)
);
wire [0:0] tree_1217;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1409 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_745),
 .b(tree_899),
 .c(tree_1217)
);
wire [0:0] tree_1218;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1410 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_655),
 .b(tree_467),
 .c(tree_1218)
);
wire [0:0] tree_1219;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1411 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_372),
 .b(tree_585),
 .c(tree_1219)
);
wire [0:0] tree_1220;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1412 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_858),
 .b(tree_552),
 .c(tree_1220)
);
wire [0:0] tree_1221;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1413 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1213),
 .b(tree_1214),
 .c(tree_1221)
);
wire [0:0] tree_1222;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1414 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1215),
 .b(tree_1216),
 .c(tree_1222)
);
wire [0:0] tree_1223;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1415 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1217),
 .b(tree_1218),
 .c(tree_1223)
);
wire [0:0] tree_1224;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1416 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1219),
 .b(tree_1220),
 .c(tree_1224)
);
wire [0:0] tree_1225;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1417 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_569),
 .b(tree_641),
 .c(tree_1225)
);
wire [0:0] tree_1226;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1418 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1221),
 .b(tree_1222),
 .c(tree_1226)
);
wire [0:0] tree_1227;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1419 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1223),
 .b(tree_1224),
 .c(tree_1227)
);
wire [0:0] tree_1228;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1420 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1225),
 .b(1'h0),
 .c(tree_1228)
);
wire [0:0] tree_1229;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1421 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1226),
 .b(tree_1227),
 .c(tree_1229)
);
wire [0:0] tree_1230;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1422 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1228),
 .b(1'h0),
 .c(tree_1230)
);
wire [0:0] tree_1231;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1423 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1229),
 .b(tree_1230),
 .c(tree_1231)
);
wire [0:0] tree_1232;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1424 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[23]),
 .b(1'h0),
 .c(tree_1232)
);
wire [0:0] tree_1233;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1425 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1232),
 .b(1'h0),
 .c(tree_1233)
);
wire [0:0] tree_1234;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1426 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1233),
 .b(tree_738),
 .c(tree_1234)
);
wire [0:0] tree_1235;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1427 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_645),
 .b(tree_665),
 .c(tree_1235)
);
wire [0:0] tree_1236;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1428 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[23]),
 .b(in[14]),
 .c(tree_1236)
);
wire [0:0] tree_1237;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1429 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[32]),
 .b(in[141]),
 .c(tree_1237)
);
wire [0:0] tree_1238;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1430 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1236),
 .b(tree_1237),
 .c(tree_1238)
);
wire [0:0] tree_1239;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1431 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_189),
 .b(tree_77),
 .c(tree_1239)
);
wire [0:0] tree_1240;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1432 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_193),
 .b(tree_376),
 .c(tree_1240)
);
wire [0:0] tree_1241;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1433 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_234),
 .b(tree_49),
 .c(tree_1241)
);
wire [0:0] tree_1242;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1434 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_117),
 .b(tree_124),
 .c(tree_1242)
);
wire [0:0] tree_1243;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1435 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_489),
 .b(tree_56),
 .c(tree_1243)
);
wire [0:0] tree_1244;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1436 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_416),
 .b(1'h0),
 .c(tree_1244)
);
wire [0:0] tree_1245;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1437 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1238),
 .b(tree_1239),
 .c(tree_1245)
);
wire [0:0] tree_1246;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1438 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1241),
 .b(tree_1240),
 .c(tree_1246)
);
wire [0:0] tree_1247;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1439 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1243),
 .b(tree_1242),
 .c(tree_1247)
);
wire [0:0] tree_1248;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1440 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1244),
 .b(tree_731),
 .c(tree_1248)
);
wire [0:0] tree_1249;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1441 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_450),
 .b(tree_998),
 .c(tree_1249)
);
wire [0:0] tree_1250;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1442 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_715),
 .b(tree_506),
 .c(tree_1250)
);
wire [0:0] tree_1251;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1443 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_549),
 .b(tree_372),
 .c(tree_1251)
);
wire [0:0] tree_1252;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1444 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_672),
 .b(tree_670),
 .c(tree_1252)
);
wire [0:0] tree_1253;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1445 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_591),
 .b(tree_316),
 .c(tree_1253)
);
wire [0:0] tree_1254;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1446 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_496),
 .b(tree_661),
 .c(tree_1254)
);
wire [0:0] tree_1255;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1447 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1245),
 .b(tree_1246),
 .c(tree_1255)
);
wire [0:0] tree_1256;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1448 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1247),
 .b(tree_1248),
 .c(tree_1256)
);
wire [0:0] tree_1257;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1449 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1249),
 .b(tree_1250),
 .c(tree_1257)
);
wire [0:0] tree_1258;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1450 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1251),
 .b(tree_1252),
 .c(tree_1258)
);
wire [0:0] tree_1259;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1451 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1253),
 .b(tree_1254),
 .c(tree_1259)
);
wire [0:0] tree_1260;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1452 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_839),
 .b(tree_675),
 .c(tree_1260)
);
wire [0:0] tree_1261;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1453 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_972),
 .b(1'h0),
 .c(tree_1261)
);
wire [0:0] tree_1262;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1454 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1255),
 .b(tree_1256),
 .c(tree_1262)
);
wire [0:0] tree_1263;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1455 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1257),
 .b(tree_1258),
 .c(tree_1263)
);
wire [0:0] tree_1264;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1456 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1259),
 .b(tree_1260),
 .c(tree_1264)
);
wire [0:0] tree_1265;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1457 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1261),
 .b(1'h0),
 .c(tree_1265)
);
wire [0:0] tree_1266;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1458 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1262),
 .b(tree_1263),
 .c(tree_1266)
);
wire [0:0] tree_1267;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1459 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1264),
 .b(tree_1265),
 .c(tree_1267)
);
wire [0:0] tree_1268;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1460 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1266),
 .b(tree_1267),
 .c(tree_1268)
);
wire [0:0] tree_1269;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1461 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_156),
 .b(1'h0),
 .c(tree_1269)
);
wire [0:0] tree_1270;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1462 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1269),
 .b(tree_677),
 .c(tree_1270)
);
wire [0:0] tree_1271;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1463 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_544),
 .b(1'h0),
 .c(tree_1271)
);
wire [0:0] tree_1272;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1464 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1271),
 .b(tree_680),
 .c(tree_1272)
);
wire [0:0] tree_1273;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1465 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[157]),
 .b(1'h0),
 .c(tree_1273)
);
wire [0:0] tree_1274;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1466 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1273),
 .b(tree_173),
 .c(tree_1274)
);
wire [0:0] tree_1275;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1467 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_335),
 .b(tree_71),
 .c(tree_1275)
);
wire [0:0] tree_1276;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1468 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_132),
 .b(tree_162),
 .c(tree_1276)
);
wire [0:0] tree_1277;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1469 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_125),
 .b(tree_222),
 .c(tree_1277)
);
wire [0:0] tree_1278;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1470 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_532),
 .b(1'h0),
 .c(tree_1278)
);
wire [0:0] tree_1279;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1471 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1275),
 .b(tree_1274),
 .c(tree_1279)
);
wire [0:0] tree_1280;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1472 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1277),
 .b(tree_1276),
 .c(tree_1280)
);
wire [0:0] tree_1281;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1473 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1278),
 .b(tree_766),
 .c(tree_1281)
);
wire [0:0] tree_1282;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1474 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_895),
 .b(tree_501),
 .c(tree_1282)
);
wire [0:0] tree_1283;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1475 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_636),
 .b(tree_802),
 .c(tree_1283)
);
wire [0:0] tree_1284;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1476 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_953),
 .b(tree_681),
 .c(tree_1284)
);
wire [0:0] tree_1285;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1477 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_656),
 .b(tree_519),
 .c(tree_1285)
);
wire [0:0] tree_1286;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1478 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_492),
 .b(tree_1031),
 .c(tree_1286)
);
wire [0:0] tree_1287;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1479 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1279),
 .b(tree_1280),
 .c(tree_1287)
);
wire [0:0] tree_1288;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1480 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1281),
 .b(tree_1282),
 .c(tree_1288)
);
wire [0:0] tree_1289;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1481 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1283),
 .b(tree_1284),
 .c(tree_1289)
);
wire [0:0] tree_1290;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1482 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1285),
 .b(tree_1286),
 .c(tree_1290)
);
wire [0:0] tree_1291;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1483 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_922),
 .b(tree_964),
 .c(tree_1291)
);
wire [0:0] tree_1292;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1484 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1287),
 .b(tree_1288),
 .c(tree_1292)
);
wire [0:0] tree_1293;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1485 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1289),
 .b(tree_1290),
 .c(tree_1293)
);
wire [0:0] tree_1294;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1486 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1291),
 .b(1'h0),
 .c(tree_1294)
);
wire [0:0] tree_1295;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1487 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1292),
 .b(tree_1293),
 .c(tree_1295)
);
wire [0:0] tree_1296;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1488 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1294),
 .b(1'h0),
 .c(tree_1296)
);
wire [0:0] tree_1297;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1489 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1295),
 .b(tree_1296),
 .c(tree_1297)
);
wire [0:0] tree_1298;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1490 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_685),
 .b(1'h0),
 .c(tree_1298)
);
wire [0:0] tree_1299;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1491 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_578),
 .b(tree_1298),
 .c(tree_1299)
);
wire [0:0] tree_1300;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1492 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_588),
 .b(1'h0),
 .c(tree_1300)
);
wire [0:0] tree_1301;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1493 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1300),
 .b(tree_944),
 .c(tree_1301)
);
wire [0:0] tree_1302;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1494 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_663),
 .b(tree_688),
 .c(tree_1302)
);
wire [0:0] tree_1303;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1495 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[29]),
 .b(in[54]),
 .c(tree_1303)
);
wire [0:0] tree_1304;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1496 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[58]),
 .b(in[170]),
 .c(tree_1304)
);
wire [0:0] tree_1305;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1497 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[178]),
 .b(1'h0),
 .c(tree_1305)
);
wire [0:0] tree_1306;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1498 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1304),
 .b(tree_1303),
 .c(tree_1306)
);
wire [0:0] tree_1307;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1499 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1305),
 .b(tree_181),
 .c(tree_1307)
);
wire [0:0] tree_1308;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1500 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_146),
 .b(tree_460),
 .c(tree_1308)
);
wire [0:0] tree_1309;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1501 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_36),
 .b(tree_57),
 .c(tree_1309)
);
wire [0:0] tree_1310;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1502 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_404),
 .b(tree_502),
 .c(tree_1310)
);
wire [0:0] tree_1311;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1503 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_579),
 .b(1'h0),
 .c(tree_1311)
);
wire [0:0] tree_1312;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1504 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1306),
 .b(tree_1307),
 .c(tree_1312)
);
wire [0:0] tree_1313;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1505 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1308),
 .b(tree_1309),
 .c(tree_1313)
);
wire [0:0] tree_1314;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1506 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1310),
 .b(tree_1311),
 .c(tree_1314)
);
wire [0:0] tree_1315;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1507 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_863),
 .b(tree_425),
 .c(tree_1315)
);
wire [0:0] tree_1316;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1508 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_436),
 .b(tree_998),
 .c(tree_1316)
);
wire [0:0] tree_1317;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1509 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_428),
 .b(tree_683),
 .c(tree_1317)
);
wire [0:0] tree_1318;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1510 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_531),
 .b(tree_1028),
 .c(tree_1318)
);
wire [0:0] tree_1319;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1511 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1104),
 .b(1'h0),
 .c(tree_1319)
);
wire [0:0] tree_1320;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1512 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1312),
 .b(tree_1313),
 .c(tree_1320)
);
wire [0:0] tree_1321;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1513 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1314),
 .b(tree_1315),
 .c(tree_1321)
);
wire [0:0] tree_1322;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1514 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1316),
 .b(tree_1317),
 .c(tree_1322)
);
wire [0:0] tree_1323;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1515 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1318),
 .b(tree_1319),
 .c(tree_1323)
);
wire [0:0] tree_1324;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1516 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1302),
 .b(1'h0),
 .c(tree_1324)
);
wire [0:0] tree_1325;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1517 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1320),
 .b(tree_1321),
 .c(tree_1325)
);
wire [0:0] tree_1326;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1518 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1322),
 .b(tree_1323),
 .c(tree_1326)
);
wire [0:0] tree_1327;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1519 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1324),
 .b(tree_1034),
 .c(tree_1327)
);
wire [0:0] tree_1328;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1520 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1325),
 .b(tree_1326),
 .c(tree_1328)
);
wire [0:0] tree_1329;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1521 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1327),
 .b(1'h0),
 .c(tree_1329)
);
wire [0:0] tree_1330;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1522 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1328),
 .b(tree_1329),
 .c(tree_1330)
);
wire [0:0] tree_1331;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1523 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_915),
 .b(tree_758),
 .c(tree_1331)
);
wire [0:0] tree_1332;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1524 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[23]),
 .b(in[121]),
 .c(tree_1332)
);
wire [0:0] tree_1333;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1525 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[165]),
 .b(in[175]),
 .c(tree_1333)
);
wire [0:0] tree_1334;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1526 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1332),
 .b(tree_1333),
 .c(tree_1334)
);
wire [0:0] tree_1335;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1527 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_86),
 .b(tree_96),
 .c(tree_1335)
);
wire [0:0] tree_1336;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1528 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_25),
 .b(tree_194),
 .c(tree_1336)
);
wire [0:0] tree_1337;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1529 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_152),
 .b(tree_122),
 .c(tree_1337)
);
wire [0:0] tree_1338;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1530 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_392),
 .b(tree_126),
 .c(tree_1338)
);
wire [0:0] tree_1339;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1531 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_161),
 .b(tree_550),
 .c(tree_1339)
);
wire [0:0] tree_1340;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1532 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_689),
 .b(tree_566),
 .c(tree_1340)
);
wire [0:0] tree_1341;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1533 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_476),
 .b(1'h0),
 .c(tree_1341)
);
wire [0:0] tree_1342;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1534 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1334),
 .b(tree_1335),
 .c(tree_1342)
);
wire [0:0] tree_1343;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1535 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1336),
 .b(tree_1337),
 .c(tree_1343)
);
wire [0:0] tree_1344;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1536 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1338),
 .b(tree_1339),
 .c(tree_1344)
);
wire [0:0] tree_1345;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1537 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1340),
 .b(tree_1341),
 .c(tree_1345)
);
wire [0:0] tree_1346;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1538 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_438),
 .b(tree_715),
 .c(tree_1346)
);
wire [0:0] tree_1347;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1539 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_563),
 .b(tree_197),
 .c(tree_1347)
);
wire [0:0] tree_1348;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1540 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_892),
 .b(tree_365),
 .c(tree_1348)
);
wire [0:0] tree_1349;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1541 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1342),
 .b(tree_1343),
 .c(tree_1349)
);
wire [0:0] tree_1350;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1542 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1344),
 .b(tree_1345),
 .c(tree_1350)
);
wire [0:0] tree_1351;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1543 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1347),
 .b(tree_1346),
 .c(tree_1351)
);
wire [0:0] tree_1352;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1544 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1348),
 .b(tree_1201),
 .c(tree_1352)
);
wire [0:0] tree_1353;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1545 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1112),
 .b(tree_979),
 .c(tree_1353)
);
wire [0:0] tree_1354;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1546 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1301),
 .b(1'h0),
 .c(tree_1354)
);
wire [0:0] tree_1355;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1547 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1349),
 .b(tree_1350),
 .c(tree_1355)
);
wire [0:0] tree_1356;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1548 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1351),
 .b(tree_1352),
 .c(tree_1356)
);
wire [0:0] tree_1357;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1549 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1353),
 .b(tree_1354),
 .c(tree_1357)
);
wire [0:0] tree_1358;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1550 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1355),
 .b(tree_1356),
 .c(tree_1358)
);
wire [0:0] tree_1359;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1551 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1357),
 .b(1'h0),
 .c(tree_1359)
);
wire [0:0] tree_1360;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1552 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1358),
 .b(tree_1359),
 .c(tree_1360)
);
wire [0:0] tree_1361;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1553 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[3]),
 .b(in[25]),
 .c(tree_1361)
);
wire [0:0] tree_1362;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1554 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1361),
 .b(tree_35),
 .c(tree_1362)
);
wire [0:0] tree_1363;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1555 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_285),
 .b(tree_249),
 .c(tree_1363)
);
wire [0:0] tree_1364;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1556 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_182),
 .b(tree_195),
 .c(tree_1364)
);
wire [0:0] tree_1365;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1557 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_361),
 .b(tree_117),
 .c(tree_1365)
);
wire [0:0] tree_1366;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1558 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_302),
 .b(tree_57),
 .c(tree_1366)
);
wire [0:0] tree_1367;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1559 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_150),
 .b(1'h0),
 .c(tree_1367)
);
wire [0:0] tree_1368;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1560 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1362),
 .b(tree_1363),
 .c(tree_1368)
);
wire [0:0] tree_1369;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1561 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1364),
 .b(tree_1365),
 .c(tree_1369)
);
wire [0:0] tree_1370;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1562 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1366),
 .b(tree_1367),
 .c(tree_1370)
);
wire [0:0] tree_1371;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1563 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_576),
 .b(tree_889),
 .c(tree_1371)
);
wire [0:0] tree_1372;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1564 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_238),
 .b(tree_444),
 .c(tree_1372)
);
wire [0:0] tree_1373;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1565 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_670),
 .b(tree_357),
 .c(tree_1373)
);
wire [0:0] tree_1374;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1566 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_651),
 .b(tree_856),
 .c(tree_1374)
);
wire [0:0] tree_1375;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1567 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1042),
 .b(tree_648),
 .c(tree_1375)
);
wire [0:0] tree_1376;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1568 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_464),
 .b(1'h0),
 .c(tree_1376)
);
wire [0:0] tree_1377;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1569 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1369),
 .b(tree_1368),
 .c(tree_1377)
);
wire [0:0] tree_1378;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1570 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1370),
 .b(tree_1371),
 .c(tree_1378)
);
wire [0:0] tree_1379;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1571 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1373),
 .b(tree_1372),
 .c(tree_1379)
);
wire [0:0] tree_1380;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1572 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1374),
 .b(tree_1375),
 .c(tree_1380)
);
wire [0:0] tree_1381;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1573 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1376),
 .b(tree_1113),
 .c(tree_1381)
);
wire [0:0] tree_1382;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1574 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1037),
 .b(1'h0),
 .c(tree_1382)
);
wire [0:0] tree_1383;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1575 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1377),
 .b(tree_1378),
 .c(tree_1383)
);
wire [0:0] tree_1384;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1576 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1379),
 .b(tree_1380),
 .c(tree_1384)
);
wire [0:0] tree_1385;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1577 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1381),
 .b(tree_1382),
 .c(tree_1385)
);
wire [0:0] tree_1386;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1578 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1383),
 .b(tree_1384),
 .c(tree_1386)
);
wire [0:0] tree_1387;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1579 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1385),
 .b(1'h0),
 .c(tree_1387)
);
wire [0:0] tree_1388;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1580 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1386),
 .b(tree_1387),
 .c(tree_1388)
);
wire [0:0] tree_1389;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1581 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[58]),
 .b(in[77]),
 .c(tree_1389)
);
wire [0:0] tree_1390;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1582 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_73),
 .b(tree_1389),
 .c(tree_1390)
);
wire [0:0] tree_1391;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1583 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_105),
 .b(tree_157),
 .c(tree_1391)
);
wire [0:0] tree_1392;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1584 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_117),
 .b(tree_277),
 .c(tree_1392)
);
wire [0:0] tree_1393;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1585 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_470),
 .b(tree_368),
 .c(tree_1393)
);
wire [0:0] tree_1394;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1586 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_356),
 .b(tree_31),
 .c(tree_1394)
);
wire [0:0] tree_1395;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1587 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_689),
 .b(tree_690),
 .c(tree_1395)
);
wire [0:0] tree_1396;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1588 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_518),
 .b(1'h0),
 .c(tree_1396)
);
wire [0:0] tree_1397;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1589 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1390),
 .b(tree_1391),
 .c(tree_1397)
);
wire [0:0] tree_1398;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1590 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1392),
 .b(tree_1393),
 .c(tree_1398)
);
wire [0:0] tree_1399;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1591 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1394),
 .b(tree_1395),
 .c(tree_1399)
);
wire [0:0] tree_1400;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1592 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1396),
 .b(tree_612),
 .c(tree_1400)
);
wire [0:0] tree_1401;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1593 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_436),
 .b(tree_598),
 .c(tree_1401)
);
wire [0:0] tree_1402;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1594 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_613),
 .b(tree_536),
 .c(tree_1402)
);
wire [0:0] tree_1403;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1595 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_554),
 .b(tree_857),
 .c(tree_1403)
);
wire [0:0] tree_1404;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1596 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_610),
 .b(1'h0),
 .c(tree_1404)
);
wire [0:0] tree_1405;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1597 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1397),
 .b(tree_1398),
 .c(tree_1405)
);
wire [0:0] tree_1406;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1598 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1399),
 .b(tree_1400),
 .c(tree_1406)
);
wire [0:0] tree_1407;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1599 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1401),
 .b(tree_1402),
 .c(tree_1407)
);
wire [0:0] tree_1408;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1600 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1403),
 .b(tree_1404),
 .c(tree_1408)
);
wire [0:0] tree_1409;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1601 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_771),
 .b(tree_884),
 .c(tree_1409)
);
wire [0:0] tree_1410;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1602 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_980),
 .b(tree_1299),
 .c(tree_1410)
);
wire [0:0] tree_1411;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1603 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1272),
 .b(1'h0),
 .c(tree_1411)
);
wire [0:0] tree_1412;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1604 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1405),
 .b(tree_1406),
 .c(tree_1412)
);
wire [0:0] tree_1413;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1605 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1407),
 .b(tree_1408),
 .c(tree_1413)
);
wire [0:0] tree_1414;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1606 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1409),
 .b(tree_1410),
 .c(tree_1414)
);
wire [0:0] tree_1415;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1607 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1411),
 .b(1'h0),
 .c(tree_1415)
);
wire [0:0] tree_1416;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1608 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1412),
 .b(tree_1413),
 .c(tree_1416)
);
wire [0:0] tree_1417;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1609 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1414),
 .b(tree_1415),
 .c(tree_1417)
);
wire [0:0] tree_1418;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1610 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1416),
 .b(tree_1417),
 .c(tree_1418)
);
wire [0:0] tree_1419;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1611 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[128]),
 .b(in[134]),
 .c(tree_1419)
);
wire [0:0] tree_1420;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1612 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[165]),
 .b(1'h0),
 .c(tree_1420)
);
wire [0:0] tree_1421;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1613 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1419),
 .b(tree_1420),
 .c(tree_1421)
);
wire [0:0] tree_1422;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1614 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_400),
 .b(tree_583),
 .c(tree_1422)
);
wire [0:0] tree_1423;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1615 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_184),
 .b(tree_596),
 .c(tree_1423)
);
wire [0:0] tree_1424;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1616 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_684),
 .b(tree_614),
 .c(tree_1424)
);
wire [0:0] tree_1425;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1617 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_653),
 .b(tree_690),
 .c(tree_1425)
);
wire [0:0] tree_1426;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1618 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1421),
 .b(tree_1422),
 .c(tree_1426)
);
wire [0:0] tree_1427;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1619 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1423),
 .b(tree_1424),
 .c(tree_1427)
);
wire [0:0] tree_1428;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1620 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_304),
 .b(tree_1425),
 .c(tree_1428)
);
wire [0:0] tree_1429;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1621 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_430),
 .b(tree_549),
 .c(tree_1429)
);
wire [0:0] tree_1430;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1622 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_951),
 .b(tree_809),
 .c(tree_1430)
);
wire [0:0] tree_1431;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1623 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_204),
 .b(tree_861),
 .c(tree_1431)
);
wire [0:0] tree_1432;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1624 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1426),
 .b(tree_1427),
 .c(tree_1432)
);
wire [0:0] tree_1433;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1625 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1428),
 .b(tree_1429),
 .c(tree_1433)
);
wire [0:0] tree_1434;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1626 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1431),
 .b(tree_1430),
 .c(tree_1434)
);
wire [0:0] tree_1435;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1627 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1331),
 .b(tree_482),
 .c(tree_1435)
);
wire [0:0] tree_1436;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1628 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1235),
 .b(tree_1270),
 .c(tree_1436)
);
wire [0:0] tree_1437;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1629 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_938),
 .b(1'h0),
 .c(tree_1437)
);
wire [0:0] tree_1438;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1630 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1432),
 .b(tree_1433),
 .c(tree_1438)
);
wire [0:0] tree_1439;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1631 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1434),
 .b(tree_1435),
 .c(tree_1439)
);
wire [0:0] tree_1440;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1632 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1436),
 .b(tree_1437),
 .c(tree_1440)
);
wire [0:0] tree_1441;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1633 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1438),
 .b(tree_1439),
 .c(tree_1441)
);
wire [0:0] tree_1442;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1634 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1440),
 .b(1'h0),
 .c(tree_1442)
);
wire [0:0] tree_1443;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1635 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1441),
 .b(tree_1442),
 .c(tree_1443)
);
wire [0:0] tree_1444;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1636 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_22),
 .b(1'h0),
 .c(tree_1444)
);
wire [0:0] tree_1445;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1637 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1444),
 .b(tree_704),
 .c(tree_1445)
);
wire [0:0] tree_1446;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1638 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_25),
 .b(1'h0),
 .c(tree_1446)
);
wire [0:0] tree_1447;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1639 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1446),
 .b(tree_706),
 .c(tree_1447)
);
wire [0:0] tree_1448;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1640 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_27),
 .b(1'h0),
 .c(tree_1448)
);
wire [0:0] tree_1449;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1641 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1448),
 .b(tree_707),
 .c(tree_1449)
);
wire [0:0] tree_1450;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1642 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_31),
 .b(1'h0),
 .c(tree_1450)
);
wire [0:0] tree_1451;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1643 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1450),
 .b(tree_709),
 .c(tree_1451)
);
wire [0:0] tree_1452;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1644 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_50),
 .b(1'h0),
 .c(tree_1452)
);
wire [0:0] tree_1453;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1645 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1452),
 .b(tree_729),
 .c(tree_1453)
);
wire [0:0] tree_1454;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1646 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_52),
 .b(1'h0),
 .c(tree_1454)
);
wire [0:0] tree_1455;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1647 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1454),
 .b(tree_731),
 .c(tree_1455)
);
wire [0:0] tree_1456;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1648 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_54),
 .b(1'h0),
 .c(tree_1456)
);
wire [0:0] tree_1457;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1649 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1456),
 .b(tree_733),
 .c(tree_1457)
);
wire [0:0] tree_1458;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1650 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[109]),
 .b(1'h0),
 .c(tree_1458)
);
wire [0:0] tree_1459;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1651 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1458),
 .b(1'h0),
 .c(tree_1459)
);
wire [0:0] tree_1460;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1652 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1459),
 .b(tree_743),
 .c(tree_1460)
);
wire [0:0] tree_1461;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1653 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_749),
 .b(tree_751),
 .c(tree_1461)
);
wire [0:0] tree_1462;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1654 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_764),
 .b(tree_766),
 .c(tree_1462)
);
wire [0:0] tree_1463;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1655 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_777),
 .b(tree_779),
 .c(tree_1463)
);
wire [0:0] tree_1464;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1656 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[53]),
 .b(in[5]),
 .c(tree_1464)
);
wire [0:0] tree_1465;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1657 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[72]),
 .b(in[109]),
 .c(tree_1465)
);
wire [0:0] tree_1466;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1658 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1464),
 .b(tree_1465),
 .c(tree_1466)
);
wire [0:0] tree_1467;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1659 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_76),
 .b(tree_35),
 .c(tree_1467)
);
wire [0:0] tree_1468;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1660 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_103),
 .b(tree_104),
 .c(tree_1468)
);
wire [0:0] tree_1469;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1661 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_105),
 .b(tree_106),
 .c(tree_1469)
);
wire [0:0] tree_1470;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1662 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_33),
 .b(tree_64),
 .c(tree_1470)
);
wire [0:0] tree_1471;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1663 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_113),
 .b(tree_112),
 .c(tree_1471)
);
wire [0:0] tree_1472;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1664 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_114),
 .b(1'h0),
 .c(tree_1472)
);
wire [0:0] tree_1473;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1665 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1466),
 .b(tree_1467),
 .c(tree_1473)
);
wire [0:0] tree_1474;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1666 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1469),
 .b(tree_1468),
 .c(tree_1474)
);
wire [0:0] tree_1475;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1667 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1470),
 .b(tree_1471),
 .c(tree_1475)
);
wire [0:0] tree_1476;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1668 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_782),
 .b(tree_1472),
 .c(tree_1476)
);
wire [0:0] tree_1477;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1669 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_784),
 .b(tree_110),
 .c(tree_1477)
);
wire [0:0] tree_1478;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1670 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_790),
 .b(tree_786),
 .c(tree_1478)
);
wire [0:0] tree_1479;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1671 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_791),
 .b(tree_792),
 .c(tree_1479)
);
wire [0:0] tree_1480;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1672 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1473),
 .b(tree_1474),
 .c(tree_1480)
);
wire [0:0] tree_1481;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1673 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1475),
 .b(tree_1476),
 .c(tree_1481)
);
wire [0:0] tree_1482;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1674 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1477),
 .b(tree_1478),
 .c(tree_1482)
);
wire [0:0] tree_1483;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1675 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1479),
 .b(tree_789),
 .c(tree_1483)
);
wire [0:0] tree_1484;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1676 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_794),
 .b(tree_1449),
 .c(tree_1484)
);
wire [0:0] tree_1485;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1677 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1480),
 .b(tree_1481),
 .c(tree_1485)
);
wire [0:0] tree_1486;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1678 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1482),
 .b(tree_1483),
 .c(tree_1486)
);
wire [0:0] tree_1487;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1679 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1484),
 .b(1'h0),
 .c(tree_1487)
);
wire [0:0] tree_1488;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1680 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1485),
 .b(tree_1486),
 .c(tree_1488)
);
wire [0:0] tree_1489;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1681 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1487),
 .b(1'h0),
 .c(tree_1489)
);
wire [0:0] tree_1490;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1682 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1488),
 .b(tree_1489),
 .c(tree_1490)
);
wire [0:0] tree_1491;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1683 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_146),
 .b(1'h0),
 .c(tree_1491)
);
wire [0:0] tree_1492;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1684 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1491),
 .b(tree_811),
 .c(tree_1492)
);
wire [0:0] tree_1493;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1685 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_829),
 .b(tree_830),
 .c(tree_1493)
);
wire [0:0] tree_1494;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1686 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[110]),
 .b(1'h0),
 .c(tree_1494)
);
wire [0:0] tree_1495;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1687 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1494),
 .b(1'h0),
 .c(tree_1495)
);
wire [0:0] tree_1496;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1688 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1495),
 .b(tree_832),
 .c(tree_1496)
);
wire [0:0] tree_1497;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1689 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_169),
 .b(1'h0),
 .c(tree_1497)
);
wire [0:0] tree_1498;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1690 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1497),
 .b(1'h0),
 .c(tree_1498)
);
wire [0:0] tree_1499;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1691 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1498),
 .b(tree_834),
 .c(tree_1499)
);
wire [0:0] tree_1500;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1692 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_181),
 .b(1'h0),
 .c(tree_1500)
);
wire [0:0] tree_1501;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1693 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1500),
 .b(tree_844),
 .c(tree_1501)
);
wire [0:0] tree_1502;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1694 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_183),
 .b(1'h0),
 .c(tree_1502)
);
wire [0:0] tree_1503;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1695 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1502),
 .b(tree_845),
 .c(tree_1503)
);
wire [0:0] tree_1504;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1696 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_188),
 .b(1'h0),
 .c(tree_1504)
);
wire [0:0] tree_1505;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1697 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1504),
 .b(tree_848),
 .c(tree_1505)
);
wire [0:0] tree_1506;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1698 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[1]),
 .b(in[26]),
 .c(tree_1506)
);
wire [0:0] tree_1507;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1699 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[143]),
 .b(1'h0),
 .c(tree_1507)
);
wire [0:0] tree_1508;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1700 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1506),
 .b(tree_1507),
 .c(tree_1508)
);
wire [0:0] tree_1509;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1701 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_173),
 .b(tree_77),
 .c(tree_1509)
);
wire [0:0] tree_1510;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1702 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_89),
 .b(tree_3),
 .c(tree_1510)
);
wire [0:0] tree_1511;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1703 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_190),
 .b(tree_158),
 .c(tree_1511)
);
wire [0:0] tree_1512;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1704 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_170),
 .b(tree_191),
 .c(tree_1512)
);
wire [0:0] tree_1513;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1705 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_155),
 .b(tree_192),
 .c(tree_1513)
);
wire [0:0] tree_1514;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1706 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_66),
 .b(1'h0),
 .c(tree_1514)
);
wire [0:0] tree_1515;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1707 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1508),
 .b(tree_1509),
 .c(tree_1515)
);
wire [0:0] tree_1516;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1708 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1511),
 .b(tree_1510),
 .c(tree_1516)
);
wire [0:0] tree_1517;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1709 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1513),
 .b(tree_1512),
 .c(tree_1517)
);
wire [0:0] tree_1518;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1710 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1514),
 .b(tree_782),
 .c(tree_1518)
);
wire [0:0] tree_1519;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1711 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_755),
 .b(tree_850),
 .c(tree_1519)
);
wire [0:0] tree_1520;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1712 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_852),
 .b(tree_853),
 .c(tree_1520)
);
wire [0:0] tree_1521;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1713 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_704),
 .b(tree_197),
 .c(tree_1521)
);
wire [0:0] tree_1522;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1714 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_855),
 .b(tree_200),
 .c(tree_1522)
);
wire [0:0] tree_1523;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1715 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_857),
 .b(tree_856),
 .c(tree_1523)
);
wire [0:0] tree_1524;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1716 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_204),
 .b(tree_858),
 .c(tree_1524)
);
wire [0:0] tree_1525;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1717 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_861),
 .b(1'h0),
 .c(tree_1525)
);
wire [0:0] tree_1526;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1718 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1515),
 .b(tree_1516),
 .c(tree_1526)
);
wire [0:0] tree_1527;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1719 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1517),
 .b(tree_1518),
 .c(tree_1527)
);
wire [0:0] tree_1528;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1720 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1519),
 .b(tree_1520),
 .c(tree_1528)
);
wire [0:0] tree_1529;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1721 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1521),
 .b(tree_1522),
 .c(tree_1529)
);
wire [0:0] tree_1530;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1722 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1523),
 .b(tree_1524),
 .c(tree_1530)
);
wire [0:0] tree_1531;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1723 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1525),
 .b(tree_860),
 .c(tree_1531)
);
wire [0:0] tree_1532;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1724 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1526),
 .b(tree_1527),
 .c(tree_1532)
);
wire [0:0] tree_1533;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1725 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1528),
 .b(tree_1529),
 .c(tree_1533)
);
wire [0:0] tree_1534;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1726 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1530),
 .b(tree_1531),
 .c(tree_1534)
);
wire [0:0] tree_1535;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1727 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1532),
 .b(tree_1533),
 .c(tree_1535)
);
wire [0:0] tree_1536;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1728 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1534),
 .b(1'h0),
 .c(tree_1536)
);
wire [0:0] tree_1537;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1729 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1535),
 .b(tree_1536),
 .c(tree_1537)
);
wire [0:0] tree_1538;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1730 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_233),
 .b(1'h0),
 .c(tree_1538)
);
wire [0:0] tree_1539;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1731 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1538),
 .b(tree_878),
 .c(tree_1539)
);
wire [0:0] tree_1540;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1732 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[71]),
 .b(in[143]),
 .c(tree_1540)
);
wire [0:0] tree_1541;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1733 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[167]),
 .b(1'h0),
 .c(tree_1541)
);
wire [0:0] tree_1542;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1734 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1541),
 .b(tree_1540),
 .c(tree_1542)
);
wire [0:0] tree_1543;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1735 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_10),
 .b(tree_16),
 .c(tree_1543)
);
wire [0:0] tree_1544;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1736 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_98),
 .b(tree_101),
 .c(tree_1544)
);
wire [0:0] tree_1545;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1737 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_234),
 .b(tree_27),
 .c(tree_1545)
);
wire [0:0] tree_1546;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1738 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_235),
 .b(tree_236),
 .c(tree_1546)
);
wire [0:0] tree_1547;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1739 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_237),
 .b(tree_239),
 .c(tree_1547)
);
wire [0:0] tree_1548;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1740 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_240),
 .b(tree_241),
 .c(tree_1548)
);
wire [0:0] tree_1549;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1741 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_244),
 .b(1'h0),
 .c(tree_1549)
);
wire [0:0] tree_1550;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1742 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1542),
 .b(tree_1543),
 .c(tree_1550)
);
wire [0:0] tree_1551;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1743 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1544),
 .b(tree_1545),
 .c(tree_1551)
);
wire [0:0] tree_1552;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1744 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1546),
 .b(tree_1547),
 .c(tree_1552)
);
wire [0:0] tree_1553;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1745 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1549),
 .b(tree_1548),
 .c(tree_1553)
);
wire [0:0] tree_1554;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1746 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_882),
 .b(tree_243),
 .c(tree_1554)
);
wire [0:0] tree_1555;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1747 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_887),
 .b(tree_246),
 .c(tree_1555)
);
wire [0:0] tree_1556;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1748 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_888),
 .b(1'h0),
 .c(tree_1556)
);
wire [0:0] tree_1557;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1749 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1550),
 .b(tree_1551),
 .c(tree_1557)
);
wire [0:0] tree_1558;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1750 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1552),
 .b(tree_1553),
 .c(tree_1558)
);
wire [0:0] tree_1559;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1751 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1554),
 .b(tree_1555),
 .c(tree_1559)
);
wire [0:0] tree_1560;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1752 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1556),
 .b(tree_881),
 .c(tree_1560)
);
wire [0:0] tree_1561;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1753 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_884),
 .b(tree_886),
 .c(tree_1561)
);
wire [0:0] tree_1562;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1754 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1557),
 .b(tree_1558),
 .c(tree_1562)
);
wire [0:0] tree_1563;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1755 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1559),
 .b(tree_1560),
 .c(tree_1563)
);
wire [0:0] tree_1564;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1756 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1561),
 .b(1'h0),
 .c(tree_1564)
);
wire [0:0] tree_1565;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1757 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1562),
 .b(tree_1563),
 .c(tree_1565)
);
wire [0:0] tree_1566;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1758 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1564),
 .b(1'h0),
 .c(tree_1566)
);
wire [0:0] tree_1567;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1759 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1565),
 .b(tree_1566),
 .c(tree_1567)
);
wire [0:0] tree_1568;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1760 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_206),
 .b(1'h0),
 .c(tree_1568)
);
wire [0:0] tree_1569;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1761 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1568),
 .b(tree_895),
 .c(tree_1569)
);
wire [0:0] tree_1570;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1762 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_282),
 .b(1'h0),
 .c(tree_1570)
);
wire [0:0] tree_1571;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1763 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1570),
 .b(1'h0),
 .c(tree_1571)
);
wire [0:0] tree_1572;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1764 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1571),
 .b(tree_913),
 .c(tree_1572)
);
wire [0:0] tree_1573;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1765 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_924),
 .b(tree_853),
 .c(tree_1573)
);
wire [0:0] tree_1574;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1766 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[102]),
 .b(in[119]),
 .c(tree_1574)
);
wire [0:0] tree_1575;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1767 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1574),
 .b(tree_173),
 .c(tree_1575)
);
wire [0:0] tree_1576;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1768 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_160),
 .b(tree_0),
 .c(tree_1576)
);
wire [0:0] tree_1577;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1769 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_100),
 .b(tree_310),
 .c(tree_1577)
);
wire [0:0] tree_1578;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1770 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_80),
 .b(tree_140),
 .c(tree_1578)
);
wire [0:0] tree_1579;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1771 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_124),
 .b(tree_36),
 .c(tree_1579)
);
wire [0:0] tree_1580;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1772 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_313),
 .b(tree_312),
 .c(tree_1580)
);
wire [0:0] tree_1581;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1773 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_320),
 .b(1'h0),
 .c(tree_1581)
);
wire [0:0] tree_1582;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1774 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1576),
 .b(tree_1575),
 .c(tree_1582)
);
wire [0:0] tree_1583;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1775 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1578),
 .b(tree_1577),
 .c(tree_1583)
);
wire [0:0] tree_1584;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1776 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1580),
 .b(tree_1579),
 .c(tree_1584)
);
wire [0:0] tree_1585;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1777 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1581),
 .b(tree_756),
 .c(tree_1585)
);
wire [0:0] tree_1586;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1778 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_784),
 .b(tree_927),
 .c(tree_1586)
);
wire [0:0] tree_1587;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1779 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_315),
 .b(tree_316),
 .c(tree_1587)
);
wire [0:0] tree_1588;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1780 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_318),
 .b(tree_929),
 .c(tree_1588)
);
wire [0:0] tree_1589;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1781 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_930),
 .b(tree_810),
 .c(tree_1589)
);
wire [0:0] tree_1590;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1782 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_931),
 .b(1'h0),
 .c(tree_1590)
);
wire [0:0] tree_1591;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1783 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1582),
 .b(tree_1583),
 .c(tree_1591)
);
wire [0:0] tree_1592;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1784 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1584),
 .b(tree_1585),
 .c(tree_1592)
);
wire [0:0] tree_1593;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1785 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1586),
 .b(tree_1587),
 .c(tree_1593)
);
wire [0:0] tree_1594;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1786 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1588),
 .b(tree_1589),
 .c(tree_1594)
);
wire [0:0] tree_1595;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1787 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1590),
 .b(tree_834),
 .c(tree_1595)
);
wire [0:0] tree_1596;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1788 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1591),
 .b(tree_1592),
 .c(tree_1596)
);
wire [0:0] tree_1597;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1789 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1593),
 .b(tree_1594),
 .c(tree_1597)
);
wire [0:0] tree_1598;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1790 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1595),
 .b(1'h0),
 .c(tree_1598)
);
wire [0:0] tree_1599;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1791 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1596),
 .b(tree_1597),
 .c(tree_1599)
);
wire [0:0] tree_1600;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1792 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1598),
 .b(1'h0),
 .c(tree_1600)
);
wire [0:0] tree_1601;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1793 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1599),
 .b(tree_1600),
 .c(tree_1601)
);
wire [0:0] tree_1602;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1794 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_940),
 .b(tree_942),
 .c(tree_1602)
);
wire [0:0] tree_1603;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1795 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[90]),
 .b(1'h0),
 .c(tree_1603)
);
wire [0:0] tree_1604;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1796 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1603),
 .b(tree_285),
 .c(tree_1604)
);
wire [0:0] tree_1605;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1797 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_252),
 .b(tree_310),
 .c(tree_1605)
);
wire [0:0] tree_1606;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1798 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_336),
 .b(tree_111),
 .c(tree_1606)
);
wire [0:0] tree_1607;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1799 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_347),
 .b(tree_338),
 .c(tree_1607)
);
wire [0:0] tree_1608;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1800 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1605),
 .b(tree_1604),
 .c(tree_1608)
);
wire [0:0] tree_1609;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1801 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1606),
 .b(tree_1607),
 .c(tree_1609)
);
wire [0:0] tree_1610;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1802 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_944),
 .b(tree_855),
 .c(tree_1610)
);
wire [0:0] tree_1611;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1803 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_946),
 .b(tree_341),
 .c(tree_1611)
);
wire [0:0] tree_1612;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1804 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_246),
 .b(tree_947),
 .c(tree_1612)
);
wire [0:0] tree_1613;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1805 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_808),
 .b(tree_741),
 .c(tree_1613)
);
wire [0:0] tree_1614;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1806 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_931),
 .b(1'h0),
 .c(tree_1614)
);
wire [0:0] tree_1615;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1807 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1608),
 .b(tree_1609),
 .c(tree_1615)
);
wire [0:0] tree_1616;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1808 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1610),
 .b(tree_1611),
 .c(tree_1616)
);
wire [0:0] tree_1617;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1809 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1612),
 .b(tree_1613),
 .c(tree_1617)
);
wire [0:0] tree_1618;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1810 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1614),
 .b(tree_948),
 .c(tree_1618)
);
wire [0:0] tree_1619;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1811 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_349),
 .b(tree_949),
 .c(tree_1619)
);
wire [0:0] tree_1620;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1812 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1615),
 .b(tree_1616),
 .c(tree_1620)
);
wire [0:0] tree_1621;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1813 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1617),
 .b(tree_1618),
 .c(tree_1621)
);
wire [0:0] tree_1622;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1814 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1619),
 .b(1'h0),
 .c(tree_1622)
);
wire [0:0] tree_1623;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1815 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1620),
 .b(tree_1621),
 .c(tree_1623)
);
wire [0:0] tree_1624;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1816 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1622),
 .b(1'h0),
 .c(tree_1624)
);
wire [0:0] tree_1625;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1817 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1623),
 .b(tree_1624),
 .c(tree_1625)
);
wire [0:0] tree_1626;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1818 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[67]),
 .b(in[14]),
 .c(tree_1626)
);
wire [0:0] tree_1627;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1819 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[79]),
 .b(in[98]),
 .c(tree_1627)
);
wire [0:0] tree_1628;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1820 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[139]),
 .b(in[186]),
 .c(tree_1628)
);
wire [0:0] tree_1629;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1821 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1626),
 .b(tree_1627),
 .c(tree_1629)
);
wire [0:0] tree_1630;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1822 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1628),
 .b(tree_245),
 .c(tree_1630)
);
wire [0:0] tree_1631;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1823 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_25),
 .b(tree_170),
 .c(tree_1631)
);
wire [0:0] tree_1632;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1824 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_147),
 .b(tree_354),
 .c(tree_1632)
);
wire [0:0] tree_1633;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1825 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_342),
 .b(tree_355),
 .c(tree_1633)
);
wire [0:0] tree_1634;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1826 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_356),
 .b(tree_359),
 .c(tree_1634)
);
wire [0:0] tree_1635;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1827 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1629),
 .b(tree_1630),
 .c(tree_1635)
);
wire [0:0] tree_1636;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1828 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1631),
 .b(tree_1632),
 .c(tree_1636)
);
wire [0:0] tree_1637;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1829 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1633),
 .b(tree_1634),
 .c(tree_1637)
);
wire [0:0] tree_1638;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1830 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_711),
 .b(tree_357),
 .c(tree_1638)
);
wire [0:0] tree_1639;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1831 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_951),
 .b(tree_315),
 .c(tree_1639)
);
wire [0:0] tree_1640;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1832 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_907),
 .b(tree_953),
 .c(tree_1640)
);
wire [0:0] tree_1641;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1833 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_791),
 .b(tree_954),
 .c(tree_1641)
);
wire [0:0] tree_1642;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1834 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_365),
 .b(1'h0),
 .c(tree_1642)
);
wire [0:0] tree_1643;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1835 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1635),
 .b(tree_1636),
 .c(tree_1643)
);
wire [0:0] tree_1644;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1836 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1637),
 .b(tree_1638),
 .c(tree_1644)
);
wire [0:0] tree_1645;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1837 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1639),
 .b(tree_1640),
 .c(tree_1645)
);
wire [0:0] tree_1646;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1838 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1641),
 .b(tree_1642),
 .c(tree_1646)
);
wire [0:0] tree_1647;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1839 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_762),
 .b(tree_957),
 .c(tree_1647)
);
wire [0:0] tree_1648;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1840 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_959),
 .b(1'h0),
 .c(tree_1648)
);
wire [0:0] tree_1649;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1841 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1643),
 .b(tree_1644),
 .c(tree_1649)
);
wire [0:0] tree_1650;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1842 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1645),
 .b(tree_1646),
 .c(tree_1650)
);
wire [0:0] tree_1651;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1843 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1647),
 .b(tree_1648),
 .c(tree_1651)
);
wire [0:0] tree_1652;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1844 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1649),
 .b(tree_1650),
 .c(tree_1652)
);
wire [0:0] tree_1653;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1845 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1651),
 .b(1'h0),
 .c(tree_1653)
);
wire [0:0] tree_1654;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1846 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1652),
 .b(tree_1653),
 .c(tree_1654)
);
wire [0:0] tree_1655;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1847 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[39]),
 .b(in[69]),
 .c(tree_1655)
);
wire [0:0] tree_1656;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1848 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[118]),
 .b(in[122]),
 .c(tree_1656)
);
wire [0:0] tree_1657;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1849 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[152]),
 .b(in[132]),
 .c(tree_1657)
);
wire [0:0] tree_1658;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1850 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[155]),
 .b(1'h0),
 .c(tree_1658)
);
wire [0:0] tree_1659;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1851 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1655),
 .b(tree_1656),
 .c(tree_1659)
);
wire [0:0] tree_1660;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1852 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1657),
 .b(tree_1658),
 .c(tree_1660)
);
wire [0:0] tree_1661;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1853 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_5),
 .b(tree_172),
 .c(tree_1661)
);
wire [0:0] tree_1662;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1854 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_367),
 .b(tree_368),
 .c(tree_1662)
);
wire [0:0] tree_1663;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1855 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_377),
 .b(1'h0),
 .c(tree_1663)
);
wire [0:0] tree_1664;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1856 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1659),
 .b(tree_1660),
 .c(tree_1664)
);
wire [0:0] tree_1665;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1857 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1662),
 .b(tree_1661),
 .c(tree_1665)
);
wire [0:0] tree_1666;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1858 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1663),
 .b(tree_760),
 .c(tree_1666)
);
wire [0:0] tree_1667;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1859 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_924),
 .b(tree_357),
 .c(tree_1667)
);
wire [0:0] tree_1668;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1860 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_370),
 .b(tree_372),
 .c(tree_1668)
);
wire [0:0] tree_1669;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1861 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_961),
 .b(tree_917),
 .c(tree_1669)
);
wire [0:0] tree_1670;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1862 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_768),
 .b(tree_734),
 .c(tree_1670)
);
wire [0:0] tree_1671;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1863 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_937),
 .b(tree_962),
 .c(tree_1671)
);
wire [0:0] tree_1672;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1864 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1664),
 .b(tree_1665),
 .c(tree_1672)
);
wire [0:0] tree_1673;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1865 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1666),
 .b(tree_1667),
 .c(tree_1673)
);
wire [0:0] tree_1674;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1866 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1668),
 .b(tree_1669),
 .c(tree_1674)
);
wire [0:0] tree_1675;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1867 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1671),
 .b(tree_1670),
 .c(tree_1675)
);
wire [0:0] tree_1676;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1868 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_375),
 .b(tree_964),
 .c(tree_1676)
);
wire [0:0] tree_1677;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1869 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1672),
 .b(tree_1673),
 .c(tree_1677)
);
wire [0:0] tree_1678;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1870 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1674),
 .b(tree_1675),
 .c(tree_1678)
);
wire [0:0] tree_1679;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1871 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1676),
 .b(1'h0),
 .c(tree_1679)
);
wire [0:0] tree_1680;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1872 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1677),
 .b(tree_1678),
 .c(tree_1680)
);
wire [0:0] tree_1681;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1873 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1679),
 .b(1'h0),
 .c(tree_1681)
);
wire [0:0] tree_1682;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1874 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1680),
 .b(tree_1681),
 .c(tree_1682)
);
wire [0:0] tree_1683;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1875 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_176),
 .b(1'h0),
 .c(tree_1683)
);
wire [0:0] tree_1684;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1876 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1683),
 .b(tree_974),
 .c(tree_1684)
);
wire [0:0] tree_1685;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1877 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[30]),
 .b(in[103]),
 .c(tree_1685)
);
wire [0:0] tree_1686;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1878 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[118]),
 .b(in[120]),
 .c(tree_1686)
);
wire [0:0] tree_1687;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1879 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1685),
 .b(tree_1686),
 .c(tree_1687)
);
wire [0:0] tree_1688;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1880 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_249),
 .b(tree_126),
 .c(tree_1688)
);
wire [0:0] tree_1689;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1881 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_378),
 .b(tree_206),
 .c(tree_1689)
);
wire [0:0] tree_1690;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1882 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_401),
 .b(tree_302),
 .c(tree_1690)
);
wire [0:0] tree_1691;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1883 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_402),
 .b(tree_145),
 .c(tree_1691)
);
wire [0:0] tree_1692;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1884 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_403),
 .b(tree_404),
 .c(tree_1692)
);
wire [0:0] tree_1693;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1885 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_405),
 .b(tree_406),
 .c(tree_1693)
);
wire [0:0] tree_1694;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1886 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_63),
 .b(tree_409),
 .c(tree_1694)
);
wire [0:0] tree_1695;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1887 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_410),
 .b(1'h0),
 .c(tree_1695)
);
wire [0:0] tree_1696;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1888 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1687),
 .b(tree_1688),
 .c(tree_1696)
);
wire [0:0] tree_1697;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1889 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1689),
 .b(tree_1690),
 .c(tree_1697)
);
wire [0:0] tree_1698;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1890 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1691),
 .b(tree_1692),
 .c(tree_1698)
);
wire [0:0] tree_1699;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1891 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1693),
 .b(tree_1694),
 .c(tree_1699)
);
wire [0:0] tree_1700;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1892 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_975),
 .b(tree_1695),
 .c(tree_1700)
);
wire [0:0] tree_1701;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1893 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_255),
 .b(tree_408),
 .c(tree_1701)
);
wire [0:0] tree_1702;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1894 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_411),
 .b(tree_394),
 .c(tree_1702)
);
wire [0:0] tree_1703;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1895 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1696),
 .b(tree_1697),
 .c(tree_1703)
);
wire [0:0] tree_1704;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1896 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1698),
 .b(tree_1699),
 .c(tree_1704)
);
wire [0:0] tree_1705;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1897 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1700),
 .b(tree_1701),
 .c(tree_1705)
);
wire [0:0] tree_1706;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1898 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1702),
 .b(tree_841),
 .c(tree_1706)
);
wire [0:0] tree_1707;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1899 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_959),
 .b(tree_977),
 .c(tree_1707)
);
wire [0:0] tree_1708;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1900 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1703),
 .b(tree_1704),
 .c(tree_1708)
);
wire [0:0] tree_1709;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1901 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1705),
 .b(tree_1706),
 .c(tree_1709)
);
wire [0:0] tree_1710;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1902 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1707),
 .b(1'h0),
 .c(tree_1710)
);
wire [0:0] tree_1711;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1903 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1708),
 .b(tree_1709),
 .c(tree_1711)
);
wire [0:0] tree_1712;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1904 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1710),
 .b(1'h0),
 .c(tree_1712)
);
wire [0:0] tree_1713;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1905 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1711),
 .b(tree_1712),
 .c(tree_1713)
);
wire [0:0] tree_1714;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1906 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[27]),
 .b(in[81]),
 .c(tree_1714)
);
wire [0:0] tree_1715;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1907 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[104]),
 .b(in[161]),
 .c(tree_1715)
);
wire [0:0] tree_1716;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1908 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1714),
 .b(tree_1715),
 .c(tree_1716)
);
wire [0:0] tree_1717;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1909 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_270),
 .b(tree_249),
 .c(tree_1717)
);
wire [0:0] tree_1718;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1910 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_212),
 .b(tree_52),
 .c(tree_1718)
);
wire [0:0] tree_1719;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1911 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_412),
 .b(tree_168),
 .c(tree_1719)
);
wire [0:0] tree_1720;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1912 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_416),
 .b(tree_292),
 .c(tree_1720)
);
wire [0:0] tree_1721;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1913 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_218),
 .b(1'h0),
 .c(tree_1721)
);
wire [0:0] tree_1722;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1914 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1716),
 .b(tree_1717),
 .c(tree_1722)
);
wire [0:0] tree_1723;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1915 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1718),
 .b(tree_1719),
 .c(tree_1723)
);
wire [0:0] tree_1724;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1916 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1720),
 .b(tree_1721),
 .c(tree_1724)
);
wire [0:0] tree_1725;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1917 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_415),
 .b(tree_224),
 .c(tree_1725)
);
wire [0:0] tree_1726;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1918 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_418),
 .b(tree_287),
 .c(tree_1726)
);
wire [0:0] tree_1727;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1919 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_420),
 .b(tree_422),
 .c(tree_1727)
);
wire [0:0] tree_1728;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1920 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_423),
 .b(tree_790),
 .c(tree_1728)
);
wire [0:0] tree_1729;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1921 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_432),
 .b(tree_431),
 .c(tree_1729)
);
wire [0:0] tree_1730;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1922 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1722),
 .b(tree_1723),
 .c(tree_1730)
);
wire [0:0] tree_1731;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1923 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1724),
 .b(tree_1725),
 .c(tree_1731)
);
wire [0:0] tree_1732;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1924 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1726),
 .b(tree_1727),
 .c(tree_1732)
);
wire [0:0] tree_1733;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1925 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1728),
 .b(tree_1729),
 .c(tree_1733)
);
wire [0:0] tree_1734;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1926 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_948),
 .b(tree_979),
 .c(tree_1734)
);
wire [0:0] tree_1735;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1927 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_980),
 .b(tree_983),
 .c(tree_1735)
);
wire [0:0] tree_1736;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1928 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1730),
 .b(tree_1731),
 .c(tree_1736)
);
wire [0:0] tree_1737;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1929 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1732),
 .b(tree_1733),
 .c(tree_1737)
);
wire [0:0] tree_1738;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1930 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1734),
 .b(tree_1735),
 .c(tree_1738)
);
wire [0:0] tree_1739;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1931 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1736),
 .b(tree_1737),
 .c(tree_1739)
);
wire [0:0] tree_1740;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1932 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1738),
 .b(1'h0),
 .c(tree_1740)
);
wire [0:0] tree_1741;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1933 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1739),
 .b(tree_1740),
 .c(tree_1741)
);
wire [0:0] tree_1742;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1934 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_177),
 .b(tree_990),
 .c(tree_1742)
);
wire [0:0] tree_1743;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1935 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[37]),
 .b(in[89]),
 .c(tree_1743)
);
wire [0:0] tree_1744;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1936 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1743),
 .b(tree_9),
 .c(tree_1744)
);
wire [0:0] tree_1745;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1937 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_226),
 .b(tree_453),
 .c(tree_1745)
);
wire [0:0] tree_1746;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1938 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_457),
 .b(tree_241),
 .c(tree_1746)
);
wire [0:0] tree_1747;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1939 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1745),
 .b(tree_1744),
 .c(tree_1747)
);
wire [0:0] tree_1748;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1940 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1746),
 .b(tree_208),
 .c(tree_1748)
);
wire [0:0] tree_1749;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1941 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_897),
 .b(tree_450),
 .c(tree_1749)
);
wire [0:0] tree_1750;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1942 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_452),
 .b(tree_154),
 .c(tree_1750)
);
wire [0:0] tree_1751;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1943 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_713),
 .b(tree_817),
 .c(tree_1751)
);
wire [0:0] tree_1752;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1944 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_459),
 .b(tree_773),
 .c(tree_1752)
);
wire [0:0] tree_1753;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1945 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_740),
 .b(tree_411),
 .c(tree_1753)
);
wire [0:0] tree_1754;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1946 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_991),
 .b(tree_993),
 .c(tree_1754)
);
wire [0:0] tree_1755;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1947 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_994),
 .b(tree_464),
 .c(tree_1755)
);
wire [0:0] tree_1756;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1948 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1747),
 .b(tree_1748),
 .c(tree_1756)
);
wire [0:0] tree_1757;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1949 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1749),
 .b(tree_1750),
 .c(tree_1757)
);
wire [0:0] tree_1758;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1950 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1751),
 .b(tree_1752),
 .c(tree_1758)
);
wire [0:0] tree_1759;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1951 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1754),
 .b(tree_1753),
 .c(tree_1759)
);
wire [0:0] tree_1760;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1952 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_456),
 .b(tree_1755),
 .c(tree_1760)
);
wire [0:0] tree_1761;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1953 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_996),
 .b(tree_997),
 .c(tree_1761)
);
wire [0:0] tree_1762;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1954 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1756),
 .b(tree_1757),
 .c(tree_1762)
);
wire [0:0] tree_1763;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1955 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1758),
 .b(tree_1759),
 .c(tree_1763)
);
wire [0:0] tree_1764;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1956 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1760),
 .b(tree_1761),
 .c(tree_1764)
);
wire [0:0] tree_1765;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1957 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1762),
 .b(tree_1763),
 .c(tree_1765)
);
wire [0:0] tree_1766;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1958 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1764),
 .b(1'h0),
 .c(tree_1766)
);
wire [0:0] tree_1767;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1959 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1765),
 .b(tree_1766),
 .c(tree_1767)
);
wire [0:0] tree_1768;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1960 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[86]),
 .b(in[119]),
 .c(tree_1768)
);
wire [0:0] tree_1769;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1961 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1768),
 .b(tree_29),
 .c(tree_1769)
);
wire [0:0] tree_1770;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1962 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_108),
 .b(tree_376),
 .c(tree_1770)
);
wire [0:0] tree_1771;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1963 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_180),
 .b(tree_98),
 .c(tree_1771)
);
wire [0:0] tree_1772;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1964 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_144),
 .b(tree_279),
 .c(tree_1772)
);
wire [0:0] tree_1773;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1965 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_470),
 .b(tree_83),
 .c(tree_1773)
);
wire [0:0] tree_1774;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1966 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_457),
 .b(tree_476),
 .c(tree_1774)
);
wire [0:0] tree_1775;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1967 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1769),
 .b(tree_1770),
 .c(tree_1775)
);
wire [0:0] tree_1776;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1968 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1771),
 .b(tree_1772),
 .c(tree_1776)
);
wire [0:0] tree_1777;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1969 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1773),
 .b(tree_1774),
 .c(tree_1777)
);
wire [0:0] tree_1778;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1970 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_706),
 .b(tree_729),
 .c(tree_1778)
);
wire [0:0] tree_1779;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1971 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_998),
 .b(tree_473),
 .c(tree_1779)
);
wire [0:0] tree_1780;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1972 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_475),
 .b(tree_422),
 .c(tree_1780)
);
wire [0:0] tree_1781;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1973 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_478),
 .b(tree_480),
 .c(tree_1781)
);
wire [0:0] tree_1782;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1974 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_431),
 .b(1'h0),
 .c(tree_1782)
);
wire [0:0] tree_1783;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1975 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1775),
 .b(tree_1776),
 .c(tree_1783)
);
wire [0:0] tree_1784;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1976 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1777),
 .b(tree_1778),
 .c(tree_1784)
);
wire [0:0] tree_1785;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1977 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1779),
 .b(tree_1780),
 .c(tree_1785)
);
wire [0:0] tree_1786;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1978 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1782),
 .b(tree_1781),
 .c(tree_1786)
);
wire [0:0] tree_1787;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1979 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_482),
 .b(tree_1001),
 .c(tree_1787)
);
wire [0:0] tree_1788;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1980 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1003),
 .b(1'h0),
 .c(tree_1788)
);
wire [0:0] tree_1789;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1981 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1783),
 .b(tree_1784),
 .c(tree_1789)
);
wire [0:0] tree_1790;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1982 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1785),
 .b(tree_1786),
 .c(tree_1790)
);
wire [0:0] tree_1791;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1983 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1787),
 .b(tree_1788),
 .c(tree_1791)
);
wire [0:0] tree_1792;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1984 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1789),
 .b(tree_1790),
 .c(tree_1792)
);
wire [0:0] tree_1793;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1985 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1791),
 .b(1'h0),
 .c(tree_1793)
);
wire [0:0] tree_1794;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1986 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1792),
 .b(tree_1793),
 .c(tree_1794)
);
wire [0:0] tree_1795;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1987 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[25]),
 .b(in[68]),
 .c(tree_1795)
);
wire [0:0] tree_1796;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1988 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[126]),
 .b(in[108]),
 .c(tree_1796)
);
wire [0:0] tree_1797;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1989 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[143]),
 .b(in[184]),
 .c(tree_1797)
);
wire [0:0] tree_1798;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1990 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1795),
 .b(tree_1796),
 .c(tree_1798)
);
wire [0:0] tree_1799;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1991 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1797),
 .b(tree_97),
 .c(tree_1799)
);
wire [0:0] tree_1800;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1992 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_87),
 .b(tree_43),
 .c(tree_1800)
);
wire [0:0] tree_1801;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1993 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_74),
 .b(tree_221),
 .c(tree_1801)
);
wire [0:0] tree_1802;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1994 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_356),
 .b(1'h0),
 .c(tree_1802)
);
wire [0:0] tree_1803;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1995 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1798),
 .b(tree_1799),
 .c(tree_1803)
);
wire [0:0] tree_1804;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1996 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1800),
 .b(tree_1801),
 .c(tree_1804)
);
wire [0:0] tree_1805;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1997 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1802),
 .b(tree_927),
 .c(tree_1805)
);
wire [0:0] tree_1806;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_1998 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_273),
 .b(tree_485),
 .c(tree_1806)
);
wire [0:0] tree_1807;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_1999 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_487),
 .b(tree_341),
 .c(tree_1807)
);
wire [0:0] tree_1808;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2000 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_488),
 .b(tree_1009),
 .c(tree_1808)
);
wire [0:0] tree_1809;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2001 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_496),
 .b(tree_492),
 .c(tree_1809)
);
wire [0:0] tree_1810;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2002 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1803),
 .b(tree_1804),
 .c(tree_1810)
);
wire [0:0] tree_1811;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2003 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1805),
 .b(tree_1806),
 .c(tree_1811)
);
wire [0:0] tree_1812;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2004 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1807),
 .b(tree_1808),
 .c(tree_1812)
);
wire [0:0] tree_1813;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2005 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1809),
 .b(tree_1005),
 .c(tree_1813)
);
wire [0:0] tree_1814;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2006 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_456),
 .b(tree_1008),
 .c(tree_1814)
);
wire [0:0] tree_1815;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2007 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1011),
 .b(tree_1014),
 .c(tree_1815)
);
wire [0:0] tree_1816;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2008 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1492),
 .b(1'h0),
 .c(tree_1816)
);
wire [0:0] tree_1817;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2009 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1810),
 .b(tree_1811),
 .c(tree_1817)
);
wire [0:0] tree_1818;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2010 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1813),
 .b(tree_1812),
 .c(tree_1818)
);
wire [0:0] tree_1819;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2011 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1814),
 .b(tree_1815),
 .c(tree_1819)
);
wire [0:0] tree_1820;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2012 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1816),
 .b(1'h0),
 .c(tree_1820)
);
wire [0:0] tree_1821;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2013 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1817),
 .b(tree_1818),
 .c(tree_1821)
);
wire [0:0] tree_1822;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2014 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1819),
 .b(tree_1820),
 .c(tree_1822)
);
wire [0:0] tree_1823;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2015 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1821),
 .b(tree_1822),
 .c(tree_1823)
);
wire [0:0] tree_1824;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2016 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[82]),
 .b(in[135]),
 .c(tree_1824)
);
wire [0:0] tree_1825;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2017 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[146]),
 .b(in[136]),
 .c(tree_1825)
);
wire [0:0] tree_1826;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2018 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[149]),
 .b(in[171]),
 .c(tree_1826)
);
wire [0:0] tree_1827;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2019 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[181]),
 .b(1'h0),
 .c(tree_1827)
);
wire [0:0] tree_1828;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2020 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1824),
 .b(tree_1825),
 .c(tree_1828)
);
wire [0:0] tree_1829;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2021 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1826),
 .b(tree_1827),
 .c(tree_1829)
);
wire [0:0] tree_1830;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2022 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_395),
 .b(tree_146),
 .c(tree_1830)
);
wire [0:0] tree_1831;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2023 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_12),
 .b(tree_312),
 .c(tree_1831)
);
wire [0:0] tree_1832;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2024 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_63),
 .b(tree_508),
 .c(tree_1832)
);
wire [0:0] tree_1833;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2025 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1828),
 .b(tree_1829),
 .c(tree_1833)
);
wire [0:0] tree_1834;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2026 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1830),
 .b(tree_1831),
 .c(tree_1834)
);
wire [0:0] tree_1835;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2027 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1832),
 .b(tree_224),
 .c(tree_1835)
);
wire [0:0] tree_1836;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2028 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_501),
 .b(tree_720),
 .c(tree_1836)
);
wire [0:0] tree_1837;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2029 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_257),
 .b(tree_1015),
 .c(tree_1837)
);
wire [0:0] tree_1838;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2030 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_509),
 .b(1'h0),
 .c(tree_1838)
);
wire [0:0] tree_1839;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2031 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1833),
 .b(tree_1834),
 .c(tree_1839)
);
wire [0:0] tree_1840;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2032 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1835),
 .b(tree_1836),
 .c(tree_1840)
);
wire [0:0] tree_1841;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2033 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1837),
 .b(tree_1838),
 .c(tree_1841)
);
wire [0:0] tree_1842;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2034 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_499),
 .b(tree_1008),
 .c(tree_1842)
);
wire [0:0] tree_1843;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2035 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1017),
 .b(tree_1018),
 .c(tree_1843)
);
wire [0:0] tree_1844;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2036 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_911),
 .b(1'h0),
 .c(tree_1844)
);
wire [0:0] tree_1845;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2037 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1839),
 .b(tree_1840),
 .c(tree_1845)
);
wire [0:0] tree_1846;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2038 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1841),
 .b(tree_1842),
 .c(tree_1846)
);
wire [0:0] tree_1847;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2039 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1843),
 .b(tree_1844),
 .c(tree_1847)
);
wire [0:0] tree_1848;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2040 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1845),
 .b(tree_1846),
 .c(tree_1848)
);
wire [0:0] tree_1849;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2041 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1847),
 .b(1'h0),
 .c(tree_1849)
);
wire [0:0] tree_1850;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2042 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1848),
 .b(tree_1849),
 .c(tree_1850)
);
wire [0:0] tree_1851;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2043 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_354),
 .b(1'h0),
 .c(tree_1851)
);
wire [0:0] tree_1852;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2044 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1851),
 .b(1'h0),
 .c(tree_1852)
);
wire [0:0] tree_1853;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2045 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1852),
 .b(tree_1020),
 .c(tree_1853)
);
wire [0:0] tree_1854;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2046 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_517),
 .b(1'h0),
 .c(tree_1854)
);
wire [0:0] tree_1855;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2047 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1023),
 .b(tree_1854),
 .c(tree_1855)
);
wire [0:0] tree_1856;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2048 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[147]),
 .b(in[42]),
 .c(tree_1856)
);
wire [0:0] tree_1857;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2049 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[150]),
 .b(1'h0),
 .c(tree_1857)
);
wire [0:0] tree_1858;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2050 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1856),
 .b(tree_1857),
 .c(tree_1858)
);
wire [0:0] tree_1859;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2051 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_25),
 .b(tree_23),
 .c(tree_1859)
);
wire [0:0] tree_1860;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2052 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_462),
 .b(tree_392),
 .c(tree_1860)
);
wire [0:0] tree_1861;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2053 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_282),
 .b(tree_11),
 .c(tree_1861)
);
wire [0:0] tree_1862;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2054 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_134),
 .b(tree_19),
 .c(tree_1862)
);
wire [0:0] tree_1863;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2055 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_518),
 .b(tree_523),
 .c(tree_1863)
);
wire [0:0] tree_1864;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2056 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_508),
 .b(1'h0),
 .c(tree_1864)
);
wire [0:0] tree_1865;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2057 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1858),
 .b(tree_1859),
 .c(tree_1865)
);
wire [0:0] tree_1866;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2058 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1860),
 .b(tree_1861),
 .c(tree_1866)
);
wire [0:0] tree_1867;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2059 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1862),
 .b(tree_1863),
 .c(tree_1867)
);
wire [0:0] tree_1868;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2060 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1864),
 .b(tree_415),
 .c(tree_1868)
);
wire [0:0] tree_1869;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2061 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_782),
 .b(tree_998),
 .c(tree_1869)
);
wire [0:0] tree_1870;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2062 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_733),
 .b(tree_385),
 .c(tree_1870)
);
wire [0:0] tree_1871;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2063 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_716),
 .b(tree_823),
 .c(tree_1871)
);
wire [0:0] tree_1872;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2064 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_804),
 .b(tree_519),
 .c(tree_1872)
);
wire [0:0] tree_1873;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2065 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_522),
 .b(tree_970),
 .c(tree_1873)
);
wire [0:0] tree_1874;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2066 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1865),
 .b(tree_1866),
 .c(tree_1874)
);
wire [0:0] tree_1875;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2067 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1867),
 .b(tree_1868),
 .c(tree_1875)
);
wire [0:0] tree_1876;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2068 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1869),
 .b(tree_1870),
 .c(tree_1876)
);
wire [0:0] tree_1877;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2069 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1871),
 .b(tree_1872),
 .c(tree_1877)
);
wire [0:0] tree_1878;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2070 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1873),
 .b(tree_499),
 .c(tree_1878)
);
wire [0:0] tree_1879;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2071 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_521),
 .b(tree_1025),
 .c(tree_1879)
);
wire [0:0] tree_1880;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2072 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1874),
 .b(tree_1875),
 .c(tree_1880)
);
wire [0:0] tree_1881;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2073 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1876),
 .b(tree_1877),
 .c(tree_1881)
);
wire [0:0] tree_1882;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2074 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1878),
 .b(tree_1879),
 .c(tree_1882)
);
wire [0:0] tree_1883;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2075 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1880),
 .b(tree_1881),
 .c(tree_1883)
);
wire [0:0] tree_1884;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2076 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1882),
 .b(1'h0),
 .c(tree_1884)
);
wire [0:0] tree_1885;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2077 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1883),
 .b(tree_1884),
 .c(tree_1885)
);
wire [0:0] tree_1886;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2078 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[3]),
 .b(in[27]),
 .c(tree_1886)
);
wire [0:0] tree_1887;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2079 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[118]),
 .b(in[74]),
 .c(tree_1887)
);
wire [0:0] tree_1888;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2080 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[191]),
 .b(1'h0),
 .c(tree_1888)
);
wire [0:0] tree_1889;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2081 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1886),
 .b(tree_1887),
 .c(tree_1889)
);
wire [0:0] tree_1890;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2082 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1888),
 .b(tree_78),
 .c(tree_1890)
);
wire [0:0] tree_1891;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2083 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_160),
 .b(tree_8),
 .c(tree_1891)
);
wire [0:0] tree_1892;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2084 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_119),
 .b(tree_155),
 .c(tree_1892)
);
wire [0:0] tree_1893;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2085 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_526),
 .b(tree_387),
 .c(tree_1893)
);
wire [0:0] tree_1894;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2086 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_532),
 .b(tree_537),
 .c(tree_1894)
);
wire [0:0] tree_1895;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2087 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1889),
 .b(tree_1890),
 .c(tree_1895)
);
wire [0:0] tree_1896;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2088 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1891),
 .b(tree_1892),
 .c(tree_1896)
);
wire [0:0] tree_1897;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2089 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1894),
 .b(tree_1893),
 .c(tree_1897)
);
wire [0:0] tree_1898;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2090 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_344),
 .b(tree_289),
 .c(tree_1898)
);
wire [0:0] tree_1899;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2091 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_531),
 .b(tree_444),
 .c(tree_1899)
);
wire [0:0] tree_1900;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2092 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_389),
 .b(tree_534),
 .c(tree_1900)
);
wire [0:0] tree_1901;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2093 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1028),
 .b(tree_536),
 .c(tree_1901)
);
wire [0:0] tree_1902;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2094 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_543),
 .b(1'h0),
 .c(tree_1902)
);
wire [0:0] tree_1903;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2095 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1895),
 .b(tree_1896),
 .c(tree_1903)
);
wire [0:0] tree_1904;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2096 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1897),
 .b(tree_1898),
 .c(tree_1904)
);
wire [0:0] tree_1905;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2097 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1899),
 .b(tree_1900),
 .c(tree_1905)
);
wire [0:0] tree_1906;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2098 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1901),
 .b(tree_1902),
 .c(tree_1906)
);
wire [0:0] tree_1907;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2099 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_529),
 .b(tree_905),
 .c(tree_1907)
);
wire [0:0] tree_1908;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2100 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1027),
 .b(tree_539),
 .c(tree_1908)
);
wire [0:0] tree_1909;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2101 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_827),
 .b(1'h0),
 .c(tree_1909)
);
wire [0:0] tree_1910;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2102 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1903),
 .b(tree_1904),
 .c(tree_1910)
);
wire [0:0] tree_1911;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2103 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1905),
 .b(tree_1906),
 .c(tree_1911)
);
wire [0:0] tree_1912;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2104 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1907),
 .b(tree_1908),
 .c(tree_1912)
);
wire [0:0] tree_1913;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2105 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1909),
 .b(1'h0),
 .c(tree_1913)
);
wire [0:0] tree_1914;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2106 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1910),
 .b(tree_1911),
 .c(tree_1914)
);
wire [0:0] tree_1915;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2107 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1912),
 .b(tree_1913),
 .c(tree_1915)
);
wire [0:0] tree_1916;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2108 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1914),
 .b(tree_1915),
 .c(tree_1916)
);
wire [0:0] tree_1917;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2109 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_212),
 .b(1'h0),
 .c(tree_1917)
);
wire [0:0] tree_1918;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2110 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1917),
 .b(1'h0),
 .c(tree_1918)
);
wire [0:0] tree_1919;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2111 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1918),
 .b(tree_1462),
 .c(tree_1919)
);
wire [0:0] tree_1920;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2112 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[176]),
 .b(in[182]),
 .c(tree_1920)
);
wire [0:0] tree_1921;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2113 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_245),
 .b(tree_1920),
 .c(tree_1921)
);
wire [0:0] tree_1922;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2114 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_61),
 .b(tree_1),
 .c(tree_1922)
);
wire [0:0] tree_1923;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2115 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_185),
 .b(tree_191),
 .c(tree_1923)
);
wire [0:0] tree_1924;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2116 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_380),
 .b(tree_406),
 .c(tree_1924)
);
wire [0:0] tree_1925;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2117 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_566),
 .b(1'h0),
 .c(tree_1925)
);
wire [0:0] tree_1926;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2118 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1921),
 .b(tree_1922),
 .c(tree_1926)
);
wire [0:0] tree_1927;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2119 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1923),
 .b(tree_1924),
 .c(tree_1927)
);
wire [0:0] tree_1928;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2120 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_436),
 .b(tree_1925),
 .c(tree_1928)
);
wire [0:0] tree_1929;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2121 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_450),
 .b(tree_560),
 .c(tree_1929)
);
wire [0:0] tree_1930;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2122 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_289),
 .b(tree_927),
 .c(tree_1930)
);
wire [0:0] tree_1931;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2123 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_562),
 .b(tree_932),
 .c(tree_1931)
);
wire [0:0] tree_1932;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2124 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_563),
 .b(tree_716),
 .c(tree_1932)
);
wire [0:0] tree_1933;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2125 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_565),
 .b(tree_571),
 .c(tree_1933)
);
wire [0:0] tree_1934;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2126 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_954),
 .b(tree_887),
 .c(tree_1934)
);
wire [0:0] tree_1935;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2127 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1926),
 .b(tree_1927),
 .c(tree_1935)
);
wire [0:0] tree_1936;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2128 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1928),
 .b(tree_1929),
 .c(tree_1936)
);
wire [0:0] tree_1937;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2129 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1930),
 .b(tree_1931),
 .c(tree_1937)
);
wire [0:0] tree_1938;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2130 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1932),
 .b(tree_1933),
 .c(tree_1938)
);
wire [0:0] tree_1939;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2131 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1934),
 .b(tree_1020),
 .c(tree_1939)
);
wire [0:0] tree_1940;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2132 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_569),
 .b(tree_1011),
 .c(tree_1940)
);
wire [0:0] tree_1941;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2133 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_977),
 .b(tree_1569),
 .c(tree_1941)
);
wire [0:0] tree_1942;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2134 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1935),
 .b(tree_1936),
 .c(tree_1942)
);
wire [0:0] tree_1943;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2135 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1937),
 .b(tree_1938),
 .c(tree_1943)
);
wire [0:0] tree_1944;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2136 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1939),
 .b(tree_1940),
 .c(tree_1944)
);
wire [0:0] tree_1945;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2137 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1941),
 .b(1'h0),
 .c(tree_1945)
);
wire [0:0] tree_1946;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2138 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1942),
 .b(tree_1943),
 .c(tree_1946)
);
wire [0:0] tree_1947;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2139 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1944),
 .b(tree_1945),
 .c(tree_1947)
);
wire [0:0] tree_1948;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2140 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1946),
 .b(tree_1947),
 .c(tree_1948)
);
wire [0:0] tree_1949;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2141 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[0]),
 .b(in[52]),
 .c(tree_1949)
);
wire [0:0] tree_1950;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2142 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[172]),
 .b(in[146]),
 .c(tree_1950)
);
wire [0:0] tree_1951;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2143 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1950),
 .b(tree_1949),
 .c(tree_1951)
);
wire [0:0] tree_1952;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2144 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_270),
 .b(tree_43),
 .c(tree_1952)
);
wire [0:0] tree_1953;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2145 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_182),
 .b(tree_5),
 .c(tree_1953)
);
wire [0:0] tree_1954;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2146 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_21),
 .b(tree_572),
 .c(tree_1954)
);
wire [0:0] tree_1955;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2147 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_406),
 .b(tree_244),
 .c(tree_1955)
);
wire [0:0] tree_1956;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2148 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1951),
 .b(tree_1952),
 .c(tree_1956)
);
wire [0:0] tree_1957;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2149 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1953),
 .b(tree_1954),
 .c(tree_1957)
);
wire [0:0] tree_1958;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2150 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1955),
 .b(tree_731),
 .c(tree_1958)
);
wire [0:0] tree_1959;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2151 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_951),
 .b(tree_534),
 .c(tree_1959)
);
wire [0:0] tree_1960;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2152 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_329),
 .b(tree_574),
 .c(tree_1960)
);
wire [0:0] tree_1961;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2153 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_200),
 .b(tree_935),
 .c(tree_1961)
);
wire [0:0] tree_1962;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2154 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_993),
 .b(tree_874),
 .c(tree_1962)
);
wire [0:0] tree_1963;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2155 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1956),
 .b(tree_1957),
 .c(tree_1963)
);
wire [0:0] tree_1964;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2156 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1958),
 .b(tree_1959),
 .c(tree_1964)
);
wire [0:0] tree_1965;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2157 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1961),
 .b(tree_1960),
 .c(tree_1965)
);
wire [0:0] tree_1966;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2158 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1962),
 .b(1'h0),
 .c(tree_1966)
);
wire [0:0] tree_1967;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2159 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1963),
 .b(tree_1964),
 .c(tree_1967)
);
wire [0:0] tree_1968;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2160 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1965),
 .b(tree_1966),
 .c(tree_1968)
);
wire [0:0] tree_1969;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2161 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1853),
 .b(tree_1034),
 .c(tree_1969)
);
wire [0:0] tree_1970;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2162 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1967),
 .b(tree_1968),
 .c(tree_1970)
);
wire [0:0] tree_1971;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2163 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1969),
 .b(1'h0),
 .c(tree_1971)
);
wire [0:0] tree_1972;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2164 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1970),
 .b(tree_1971),
 .c(tree_1972)
);
wire [0:0] tree_1973;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2165 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[171]),
 .b(in[176]),
 .c(tree_1973)
);
wire [0:0] tree_1974;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2166 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[181]),
 .b(1'h0),
 .c(tree_1974)
);
wire [0:0] tree_1975;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2167 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1973),
 .b(tree_1974),
 .c(tree_1975)
);
wire [0:0] tree_1976;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2168 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_0),
 .b(tree_61),
 .c(tree_1976)
);
wire [0:0] tree_1977;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2169 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_123),
 .b(tree_16),
 .c(tree_1977)
);
wire [0:0] tree_1978;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2170 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_74),
 .b(tree_41),
 .c(tree_1978)
);
wire [0:0] tree_1979;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2171 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_405),
 .b(tree_547),
 .c(tree_1979)
);
wire [0:0] tree_1980;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2172 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_237),
 .b(tree_580),
 .c(tree_1980)
);
wire [0:0] tree_1981;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2173 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1975),
 .b(tree_1976),
 .c(tree_1981)
);
wire [0:0] tree_1982;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2174 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1977),
 .b(tree_1978),
 .c(tree_1982)
);
wire [0:0] tree_1983;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2175 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1979),
 .b(tree_1980),
 .c(tree_1983)
);
wire [0:0] tree_1984;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2176 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_515),
 .b(tree_706),
 .c(tree_1984)
);
wire [0:0] tree_1985;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2177 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_779),
 .b(tree_525),
 .c(tree_1985)
);
wire [0:0] tree_1986;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2178 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_724),
 .b(tree_818),
 .c(tree_1986)
);
wire [0:0] tree_1987;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2179 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_391),
 .b(tree_584),
 .c(tree_1987)
);
wire [0:0] tree_1988;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2180 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_991),
 .b(tree_318),
 .c(tree_1988)
);
wire [0:0] tree_1989;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2181 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1981),
 .b(tree_1982),
 .c(tree_1989)
);
wire [0:0] tree_1990;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2182 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1983),
 .b(tree_1984),
 .c(tree_1990)
);
wire [0:0] tree_1991;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2183 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1985),
 .b(tree_1986),
 .c(tree_1991)
);
wire [0:0] tree_1992;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2184 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1987),
 .b(tree_1988),
 .c(tree_1992)
);
wire [0:0] tree_1993;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2185 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_789),
 .b(tree_1037),
 .c(tree_1993)
);
wire [0:0] tree_1994;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2186 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1989),
 .b(tree_1990),
 .c(tree_1994)
);
wire [0:0] tree_1995;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2187 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1991),
 .b(tree_1992),
 .c(tree_1995)
);
wire [0:0] tree_1996;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2188 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1993),
 .b(1'h0),
 .c(tree_1996)
);
wire [0:0] tree_1997;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2189 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1994),
 .b(tree_1995),
 .c(tree_1997)
);
wire [0:0] tree_1998;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2190 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_1996),
 .b(1'h0),
 .c(tree_1998)
);
wire [0:0] tree_1999;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2191 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_1997),
 .b(tree_1998),
 .c(tree_1999)
);
wire [0:0] tree_2000;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2192 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[75]),
 .b(in[96]),
 .c(tree_2000)
);
wire [0:0] tree_2001;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2193 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[111]),
 .b(in[177]),
 .c(tree_2001)
);
wire [0:0] tree_2002;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2194 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2000),
 .b(tree_2001),
 .c(tree_2002)
);
wire [0:0] tree_2003;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2195 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_82),
 .b(tree_51),
 .c(tree_2003)
);
wire [0:0] tree_2004;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2196 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_77),
 .b(tree_252),
 .c(tree_2004)
);
wire [0:0] tree_2005;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2197 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_310),
 .b(tree_52),
 .c(tree_2005)
);
wire [0:0] tree_2006;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2198 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_361),
 .b(tree_588),
 .c(tree_2006)
);
wire [0:0] tree_2007;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2199 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_236),
 .b(tree_405),
 .c(tree_2007)
);
wire [0:0] tree_2008;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2200 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_313),
 .b(tree_259),
 .c(tree_2008)
);
wire [0:0] tree_2009;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2201 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2002),
 .b(tree_2003),
 .c(tree_2009)
);
wire [0:0] tree_2010;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2202 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2004),
 .b(tree_2005),
 .c(tree_2010)
);
wire [0:0] tree_2011;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2203 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2006),
 .b(tree_2007),
 .c(tree_2011)
);
wire [0:0] tree_2012;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2204 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2008),
 .b(tree_273),
 .c(tree_2012)
);
wire [0:0] tree_2013;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2205 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_590),
 .b(tree_562),
 .c(tree_2013)
);
wire [0:0] tree_2014;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2206 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_882),
 .b(tree_591),
 .c(tree_2014)
);
wire [0:0] tree_2015;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2207 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_592),
 .b(tree_739),
 .c(tree_2015)
);
wire [0:0] tree_2016;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2208 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_775),
 .b(1'h0),
 .c(tree_2016)
);
wire [0:0] tree_2017;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2209 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2009),
 .b(tree_2010),
 .c(tree_2017)
);
wire [0:0] tree_2018;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2210 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2011),
 .b(tree_2012),
 .c(tree_2018)
);
wire [0:0] tree_2019;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2211 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2013),
 .b(tree_2014),
 .c(tree_2019)
);
wire [0:0] tree_2020;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2212 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2015),
 .b(tree_2016),
 .c(tree_2020)
);
wire [0:0] tree_2021;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2213 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_762),
 .b(tree_499),
 .c(tree_2021)
);
wire [0:0] tree_2022;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2214 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_821),
 .b(tree_934),
 .c(tree_2022)
);
wire [0:0] tree_2023;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2215 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1742),
 .b(1'h0),
 .c(tree_2023)
);
wire [0:0] tree_2024;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2216 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2017),
 .b(tree_2018),
 .c(tree_2024)
);
wire [0:0] tree_2025;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2217 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2019),
 .b(tree_2020),
 .c(tree_2025)
);
wire [0:0] tree_2026;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2218 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2021),
 .b(tree_2022),
 .c(tree_2026)
);
wire [0:0] tree_2027;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2219 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2023),
 .b(1'h0),
 .c(tree_2027)
);
wire [0:0] tree_2028;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2220 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2024),
 .b(tree_2025),
 .c(tree_2028)
);
wire [0:0] tree_2029;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2221 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2026),
 .b(tree_2027),
 .c(tree_2029)
);
wire [0:0] tree_2030;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2222 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2028),
 .b(tree_2029),
 .c(tree_2030)
);
wire [0:0] tree_2031;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2223 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[57]),
 .b(in[17]),
 .c(tree_2031)
);
wire [0:0] tree_2032;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2224 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[117]),
 .b(1'h0),
 .c(tree_2032)
);
wire [0:0] tree_2033;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2225 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2031),
 .b(tree_2032),
 .c(tree_2033)
);
wire [0:0] tree_2034;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2226 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_201),
 .b(tree_126),
 .c(tree_2034)
);
wire [0:0] tree_2035;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2227 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_195),
 .b(tree_185),
 .c(tree_2035)
);
wire [0:0] tree_2036;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2228 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_118),
 .b(tree_462),
 .c(tree_2036)
);
wire [0:0] tree_2037;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2229 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_593),
 .b(tree_192),
 .c(tree_2037)
);
wire [0:0] tree_2038;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2230 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_594),
 .b(1'h0),
 .c(tree_2038)
);
wire [0:0] tree_2039;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2231 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2033),
 .b(tree_2034),
 .c(tree_2039)
);
wire [0:0] tree_2040;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2232 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2035),
 .b(tree_2036),
 .c(tree_2040)
);
wire [0:0] tree_2041;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2233 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2037),
 .b(tree_2038),
 .c(tree_2041)
);
wire [0:0] tree_2042;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2234 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_434),
 .b(tree_692),
 .c(tree_2042)
);
wire [0:0] tree_2043;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2235 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_546),
 .b(tree_736),
 .c(tree_2043)
);
wire [0:0] tree_2044;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2236 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_131),
 .b(tree_420),
 .c(tree_2044)
);
wire [0:0] tree_2045;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2237 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_243),
 .b(tree_774),
 .c(tree_2045)
);
wire [0:0] tree_2046;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2238 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_592),
 .b(tree_595),
 .c(tree_2046)
);
wire [0:0] tree_2047;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2239 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1041),
 .b(1'h0),
 .c(tree_2047)
);
wire [0:0] tree_2048;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2240 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2039),
 .b(tree_2040),
 .c(tree_2048)
);
wire [0:0] tree_2049;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2241 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2041),
 .b(tree_2042),
 .c(tree_2049)
);
wire [0:0] tree_2050;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2242 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2043),
 .b(tree_2044),
 .c(tree_2050)
);
wire [0:0] tree_2051;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2243 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2046),
 .b(tree_2045),
 .c(tree_2051)
);
wire [0:0] tree_2052;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2244 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2047),
 .b(tree_1040),
 .c(tree_2052)
);
wire [0:0] tree_2053;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2245 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1457),
 .b(tree_1030),
 .c(tree_2053)
);
wire [0:0] tree_2054;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2246 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2048),
 .b(tree_2049),
 .c(tree_2054)
);
wire [0:0] tree_2055;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2247 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2050),
 .b(tree_2051),
 .c(tree_2055)
);
wire [0:0] tree_2056;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2248 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2052),
 .b(tree_2053),
 .c(tree_2056)
);
wire [0:0] tree_2057;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2249 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2054),
 .b(tree_2055),
 .c(tree_2057)
);
wire [0:0] tree_2058;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2250 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2056),
 .b(1'h0),
 .c(tree_2058)
);
wire [0:0] tree_2059;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2251 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2057),
 .b(tree_2058),
 .c(tree_2059)
);
wire [0:0] tree_2060;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2252 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[53]),
 .b(in[120]),
 .c(tree_2060)
);
wire [0:0] tree_2061;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2253 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[130]),
 .b(in[152]),
 .c(tree_2061)
);
wire [0:0] tree_2062;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2254 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[163]),
 .b(in[180]),
 .c(tree_2062)
);
wire [0:0] tree_2063;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2255 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2061),
 .b(tree_2060),
 .c(tree_2063)
);
wire [0:0] tree_2064;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2256 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2062),
 .b(tree_28),
 .c(tree_2064)
);
wire [0:0] tree_2065;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2257 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_151),
 .b(tree_141),
 .c(tree_2065)
);
wire [0:0] tree_2066;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2258 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_153),
 .b(tree_198),
 .c(tree_2066)
);
wire [0:0] tree_2067;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2259 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_227),
 .b(tree_147),
 .c(tree_2067)
);
wire [0:0] tree_2068;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2260 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_136),
 .b(tree_253),
 .c(tree_2068)
);
wire [0:0] tree_2069;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2261 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_599),
 .b(tree_602),
 .c(tree_2069)
);
wire [0:0] tree_2070;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2262 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2063),
 .b(tree_2064),
 .c(tree_2070)
);
wire [0:0] tree_2071;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2263 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2065),
 .b(tree_2066),
 .c(tree_2071)
);
wire [0:0] tree_2072;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2264 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2067),
 .b(tree_2068),
 .c(tree_2072)
);
wire [0:0] tree_2073;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2265 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2069),
 .b(tree_452),
 .c(tree_2073)
);
wire [0:0] tree_2074;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2266 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_291),
 .b(tree_598),
 .c(tree_2074)
);
wire [0:0] tree_2075;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2267 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_600),
 .b(tree_220),
 .c(tree_2075)
);
wire [0:0] tree_2076;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2268 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_595),
 .b(tree_1009),
 .c(tree_2076)
);
wire [0:0] tree_2077;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2269 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1042),
 .b(1'h0),
 .c(tree_2077)
);
wire [0:0] tree_2078;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2270 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2070),
 .b(tree_2071),
 .c(tree_2078)
);
wire [0:0] tree_2079;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2271 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2072),
 .b(tree_2073),
 .c(tree_2079)
);
wire [0:0] tree_2080;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2272 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2074),
 .b(tree_2075),
 .c(tree_2080)
);
wire [0:0] tree_2081;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2273 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2076),
 .b(tree_2077),
 .c(tree_2081)
);
wire [0:0] tree_2082;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2274 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1001),
 .b(tree_902),
 .c(tree_2082)
);
wire [0:0] tree_2083;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2275 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2078),
 .b(tree_2079),
 .c(tree_2083)
);
wire [0:0] tree_2084;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2276 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2080),
 .b(tree_2081),
 .c(tree_2084)
);
wire [0:0] tree_2085;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2277 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2082),
 .b(1'h0),
 .c(tree_2085)
);
wire [0:0] tree_2086;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2278 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2083),
 .b(tree_2084),
 .c(tree_2086)
);
wire [0:0] tree_2087;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2279 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2085),
 .b(1'h0),
 .c(tree_2087)
);
wire [0:0] tree_2088;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2280 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2086),
 .b(tree_2087),
 .c(tree_2088)
);
wire [0:0] tree_2089;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2281 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[49]),
 .b(in[63]),
 .c(tree_2089)
);
wire [0:0] tree_2090;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2282 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[67]),
 .b(in[88]),
 .c(tree_2090)
);
wire [0:0] tree_2091;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2283 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2089),
 .b(tree_2090),
 .c(tree_2091)
);
wire [0:0] tree_2092;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2284 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_10),
 .b(tree_77),
 .c(tree_2092)
);
wire [0:0] tree_2093;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2285 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_164),
 .b(tree_70),
 .c(tree_2093)
);
wire [0:0] tree_2094;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2286 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_264),
 .b(tree_91),
 .c(tree_2094)
);
wire [0:0] tree_2095;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2287 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_271),
 .b(tree_470),
 .c(tree_2095)
);
wire [0:0] tree_2096;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2288 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_579),
 .b(tree_239),
 .c(tree_2096)
);
wire [0:0] tree_2097;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2289 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_621),
 .b(tree_377),
 .c(tree_2097)
);
wire [0:0] tree_2098;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2290 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2091),
 .b(tree_2092),
 .c(tree_2098)
);
wire [0:0] tree_2099;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2291 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2093),
 .b(tree_2094),
 .c(tree_2099)
);
wire [0:0] tree_2100;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2292 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2095),
 .b(tree_2096),
 .c(tree_2100)
);
wire [0:0] tree_2101;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2293 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2097),
 .b(tree_325),
 .c(tree_2101)
);
wire [0:0] tree_2102;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2294 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_620),
 .b(tree_294),
 .c(tree_2102)
);
wire [0:0] tree_2103;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2295 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_966),
 .b(tree_563),
 .c(tree_2103)
);
wire [0:0] tree_2104;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2296 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_608),
 .b(tree_613),
 .c(tree_2104)
);
wire [0:0] tree_2105;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2297 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_600),
 .b(tree_1104),
 .c(tree_2105)
);
wire [0:0] tree_2106;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2298 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_624),
 .b(tree_872),
 .c(tree_2106)
);
wire [0:0] tree_2107;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2299 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2098),
 .b(tree_2099),
 .c(tree_2107)
);
wire [0:0] tree_2108;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2300 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2100),
 .b(tree_2101),
 .c(tree_2108)
);
wire [0:0] tree_2109;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2301 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2102),
 .b(tree_2103),
 .c(tree_2109)
);
wire [0:0] tree_2110;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2302 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2104),
 .b(tree_2105),
 .c(tree_2110)
);
wire [0:0] tree_2111;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2303 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2106),
 .b(tree_997),
 .c(tree_2111)
);
wire [0:0] tree_2112;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2304 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2107),
 .b(tree_2108),
 .c(tree_2112)
);
wire [0:0] tree_2113;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2305 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2110),
 .b(tree_2109),
 .c(tree_2113)
);
wire [0:0] tree_2114;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2306 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2111),
 .b(1'h0),
 .c(tree_2114)
);
wire [0:0] tree_2115;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2307 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2112),
 .b(tree_2113),
 .c(tree_2115)
);
wire [0:0] tree_2116;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2308 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2114),
 .b(1'h0),
 .c(tree_2116)
);
wire [0:0] tree_2117;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2309 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2115),
 .b(tree_2116),
 .c(tree_2117)
);
wire [0:0] tree_2118;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2310 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[2]),
 .b(in[20]),
 .c(tree_2118)
);
wire [0:0] tree_2119;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2311 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[27]),
 .b(in[47]),
 .c(tree_2119)
);
wire [0:0] tree_2120;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2312 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[154]),
 .b(in[162]),
 .c(tree_2120)
);
wire [0:0] tree_2121;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2313 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2118),
 .b(tree_2119),
 .c(tree_2121)
);
wire [0:0] tree_2122;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2314 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2120),
 .b(tree_263),
 .c(tree_2122)
);
wire [0:0] tree_2123;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2315 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_260),
 .b(tree_40),
 .c(tree_2123)
);
wire [0:0] tree_2124;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2316 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_489),
 .b(tree_65),
 .c(tree_2124)
);
wire [0:0] tree_2125;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2317 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_347),
 .b(tree_113),
 .c(tree_2125)
);
wire [0:0] tree_2126;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2318 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2121),
 .b(tree_2122),
 .c(tree_2126)
);
wire [0:0] tree_2127;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2319 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2123),
 .b(tree_2124),
 .c(tree_2127)
);
wire [0:0] tree_2128;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2320 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2125),
 .b(tree_764),
 .c(tree_2128)
);
wire [0:0] tree_2129;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2321 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_755),
 .b(tree_696),
 .c(tree_2129)
);
wire [0:0] tree_2130;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2322 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_187),
 .b(tree_450),
 .c(tree_2130)
);
wire [0:0] tree_2131;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2323 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_268),
 .b(tree_814),
 .c(tree_2131)
);
wire [0:0] tree_2132;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2324 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_930),
 .b(1'h0),
 .c(tree_2132)
);
wire [0:0] tree_2133;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2325 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2126),
 .b(tree_2127),
 .c(tree_2133)
);
wire [0:0] tree_2134;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2326 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2128),
 .b(tree_2129),
 .c(tree_2134)
);
wire [0:0] tree_2135;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2327 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2130),
 .b(tree_2131),
 .c(tree_2135)
);
wire [0:0] tree_2136;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2328 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2132),
 .b(tree_920),
 .c(tree_2136)
);
wire [0:0] tree_2137;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2329 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1110),
 .b(tree_626),
 .c(tree_2137)
);
wire [0:0] tree_2138;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2330 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1014),
 .b(1'h0),
 .c(tree_2138)
);
wire [0:0] tree_2139;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2331 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2133),
 .b(tree_2134),
 .c(tree_2139)
);
wire [0:0] tree_2140;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2332 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2135),
 .b(tree_2136),
 .c(tree_2140)
);
wire [0:0] tree_2141;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2333 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2137),
 .b(tree_2138),
 .c(tree_2141)
);
wire [0:0] tree_2142;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2334 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1108),
 .b(1'h0),
 .c(tree_2142)
);
wire [0:0] tree_2143;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2335 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2139),
 .b(tree_2140),
 .c(tree_2143)
);
wire [0:0] tree_2144;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2336 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2141),
 .b(tree_2142),
 .c(tree_2144)
);
wire [0:0] tree_2145;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2337 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2143),
 .b(tree_2144),
 .c(tree_2145)
);
wire [0:0] tree_2146;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2338 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[96]),
 .b(in[57]),
 .c(tree_2146)
);
wire [0:0] tree_2147;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2339 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[115]),
 .b(in[100]),
 .c(tree_2147)
);
wire [0:0] tree_2148;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2340 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2146),
 .b(tree_2147),
 .c(tree_2148)
);
wire [0:0] tree_2149;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2341 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_103),
 .b(tree_88),
 .c(tree_2149)
);
wire [0:0] tree_2150;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2342 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_339),
 .b(tree_6),
 .c(tree_2150)
);
wire [0:0] tree_2151;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2343 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_337),
 .b(tree_265),
 .c(tree_2151)
);
wire [0:0] tree_2152;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2344 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_8),
 .b(tree_355),
 .c(tree_2152)
);
wire [0:0] tree_2153;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2345 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_368),
 .b(tree_114),
 .c(tree_2153)
);
wire [0:0] tree_2154;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2346 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2148),
 .b(tree_2149),
 .c(tree_2154)
);
wire [0:0] tree_2155;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2347 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2150),
 .b(tree_2151),
 .c(tree_2155)
);
wire [0:0] tree_2156;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2348 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2153),
 .b(tree_2152),
 .c(tree_2156)
);
wire [0:0] tree_2157;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2349 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_758),
 .b(tree_558),
 .c(tree_2157)
);
wire [0:0] tree_2158;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2350 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_301),
 .b(tree_582),
 .c(tree_2158)
);
wire [0:0] tree_2159;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2351 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_616),
 .b(tree_726),
 .c(tree_2159)
);
wire [0:0] tree_2160;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2352 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_624),
 .b(1'h0),
 .c(tree_2160)
);
wire [0:0] tree_2161;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2353 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2154),
 .b(tree_2155),
 .c(tree_2161)
);
wire [0:0] tree_2162;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2354 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2156),
 .b(tree_2157),
 .c(tree_2162)
);
wire [0:0] tree_2163;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2355 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2159),
 .b(tree_2158),
 .c(tree_2163)
);
wire [0:0] tree_2164;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2356 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2160),
 .b(tree_1460),
 .c(tree_2164)
);
wire [0:0] tree_2165;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2357 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_989),
 .b(tree_1112),
 .c(tree_2165)
);
wire [0:0] tree_2166;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2358 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1115),
 .b(tree_1113),
 .c(tree_2166)
);
wire [0:0] tree_2167;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2359 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1117),
 .b(1'h0),
 .c(tree_2167)
);
wire [0:0] tree_2168;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2360 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2161),
 .b(tree_2162),
 .c(tree_2168)
);
wire [0:0] tree_2169;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2361 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2163),
 .b(tree_2164),
 .c(tree_2169)
);
wire [0:0] tree_2170;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2362 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2165),
 .b(tree_2166),
 .c(tree_2170)
);
wire [0:0] tree_2171;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2363 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2167),
 .b(tree_1108),
 .c(tree_2171)
);
wire [0:0] tree_2172;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2364 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2168),
 .b(tree_2169),
 .c(tree_2172)
);
wire [0:0] tree_2173;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2365 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2170),
 .b(tree_2171),
 .c(tree_2173)
);
wire [0:0] tree_2174;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2366 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2172),
 .b(tree_2173),
 .c(tree_2174)
);
wire [0:0] tree_2175;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2367 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[81]),
 .b(in[107]),
 .c(tree_2175)
);
wire [0:0] tree_2176;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2368 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[115]),
 .b(1'h0),
 .c(tree_2176)
);
wire [0:0] tree_2177;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2369 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2175),
 .b(tree_2176),
 .c(tree_2177)
);
wire [0:0] tree_2178;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2370 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_160),
 .b(tree_310),
 .c(tree_2178)
);
wire [0:0] tree_2179;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2371 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_209),
 .b(tree_47),
 .c(tree_2179)
);
wire [0:0] tree_2180;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2372 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_652),
 .b(tree_653),
 .c(tree_2180)
);
wire [0:0] tree_2181;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2373 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2177),
 .b(tree_2178),
 .c(tree_2181)
);
wire [0:0] tree_2182;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2374 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2179),
 .b(tree_2180),
 .c(tree_2182)
);
wire [0:0] tree_2183;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2375 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_187),
 .b(tree_829),
 .c(tree_2183)
);
wire [0:0] tree_2184;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2376 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_844),
 .b(tree_217),
 .c(tree_2184)
);
wire [0:0] tree_2185;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2377 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_571),
 .b(tree_651),
 .c(tree_2185)
);
wire [0:0] tree_2186;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2378 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_968),
 .b(tree_921),
 .c(tree_2186)
);
wire [0:0] tree_2187;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2379 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_656),
 .b(1'h0),
 .c(tree_2187)
);
wire [0:0] tree_2188;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2380 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2181),
 .b(tree_2182),
 .c(tree_2188)
);
wire [0:0] tree_2189;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2381 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2183),
 .b(tree_2184),
 .c(tree_2189)
);
wire [0:0] tree_2190;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2382 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2185),
 .b(tree_2186),
 .c(tree_2190)
);
wire [0:0] tree_2191;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2383 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2187),
 .b(tree_1201),
 .c(tree_2191)
);
wire [0:0] tree_2192;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2384 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1453),
 .b(tree_521),
 .c(tree_2192)
);
wire [0:0] tree_2193;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2385 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1025),
 .b(tree_1202),
 .c(tree_2193)
);
wire [0:0] tree_2194;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2386 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2188),
 .b(tree_2189),
 .c(tree_2194)
);
wire [0:0] tree_2195;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2387 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2190),
 .b(tree_2191),
 .c(tree_2195)
);
wire [0:0] tree_2196;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2388 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2192),
 .b(tree_2193),
 .c(tree_2196)
);
wire [0:0] tree_2197;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2389 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2194),
 .b(tree_2195),
 .c(tree_2197)
);
wire [0:0] tree_2198;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2390 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2196),
 .b(1'h0),
 .c(tree_2198)
);
wire [0:0] tree_2199;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2391 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2197),
 .b(tree_2198),
 .c(tree_2199)
);
wire [0:0] tree_2200;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2392 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[3]),
 .b(in[52]),
 .c(tree_2200)
);
wire [0:0] tree_2201;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2393 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[92]),
 .b(in[84]),
 .c(tree_2201)
);
wire [0:0] tree_2202;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2394 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2200),
 .b(tree_2201),
 .c(tree_2202)
);
wire [0:0] tree_2203;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2395 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_49),
 .b(tree_383),
 .c(tree_2203)
);
wire [0:0] tree_2204;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2396 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_260),
 .b(tree_460),
 .c(tree_2204)
);
wire [0:0] tree_2205;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2397 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_652),
 .b(tree_403),
 .c(tree_2205)
);
wire [0:0] tree_2206;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2398 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_269),
 .b(1'h0),
 .c(tree_2206)
);
wire [0:0] tree_2207;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2399 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2202),
 .b(tree_2203),
 .c(tree_2207)
);
wire [0:0] tree_2208;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2400 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2204),
 .b(tree_2205),
 .c(tree_2208)
);
wire [0:0] tree_2209;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2401 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_711),
 .b(tree_2206),
 .c(tree_2209)
);
wire [0:0] tree_2210;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2402 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_284),
 .b(tree_370),
 .c(tree_2210)
);
wire [0:0] tree_2211;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2403 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_658),
 .b(tree_1036),
 .c(tree_2211)
);
wire [0:0] tree_2212;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2404 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_660),
 .b(tree_807),
 .c(tree_2212)
);
wire [0:0] tree_2213;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2405 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_661),
 .b(tree_909),
 .c(tree_2213)
);
wire [0:0] tree_2214;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2406 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_143),
 .b(tree_543),
 .c(tree_2214)
);
wire [0:0] tree_2215;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2407 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_649),
 .b(tree_873),
 .c(tree_2215)
);
wire [0:0] tree_2216;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2408 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_962),
 .b(1'h0),
 .c(tree_2216)
);
wire [0:0] tree_2217;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2409 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2207),
 .b(tree_2208),
 .c(tree_2217)
);
wire [0:0] tree_2218;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2410 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2209),
 .b(tree_2210),
 .c(tree_2218)
);
wire [0:0] tree_2219;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2411 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2211),
 .b(tree_2212),
 .c(tree_2219)
);
wire [0:0] tree_2220;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2412 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2213),
 .b(tree_2214),
 .c(tree_2220)
);
wire [0:0] tree_2221;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2413 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2215),
 .b(tree_2216),
 .c(tree_2221)
);
wire [0:0] tree_2222;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2414 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1040),
 .b(tree_1203),
 .c(tree_2222)
);
wire [0:0] tree_2223;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2415 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_349),
 .b(1'h0),
 .c(tree_2223)
);
wire [0:0] tree_2224;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2416 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2217),
 .b(tree_2218),
 .c(tree_2224)
);
wire [0:0] tree_2225;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2417 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2219),
 .b(tree_2220),
 .c(tree_2225)
);
wire [0:0] tree_2226;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2418 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2222),
 .b(tree_2221),
 .c(tree_2226)
);
wire [0:0] tree_2227;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2419 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2223),
 .b(1'h0),
 .c(tree_2227)
);
wire [0:0] tree_2228;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2420 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2224),
 .b(tree_2225),
 .c(tree_2228)
);
wire [0:0] tree_2229;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2421 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2226),
 .b(tree_2227),
 .c(tree_2229)
);
wire [0:0] tree_2230;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2422 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2228),
 .b(tree_2229),
 .c(tree_2230)
);
wire [0:0] tree_2231;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2423 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[42]),
 .b(in[90]),
 .c(tree_2231)
);
wire [0:0] tree_2232;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2424 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[109]),
 .b(in[116]),
 .c(tree_2232)
);
wire [0:0] tree_2233;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2425 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[173]),
 .b(in[137]),
 .c(tree_2233)
);
wire [0:0] tree_2234;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2426 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[185]),
 .b(1'h0),
 .c(tree_2234)
);
wire [0:0] tree_2235;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2427 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2231),
 .b(tree_2232),
 .c(tree_2235)
);
wire [0:0] tree_2236;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2428 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2233),
 .b(tree_2234),
 .c(tree_2236)
);
wire [0:0] tree_2237;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2429 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_84),
 .b(tree_360),
 .c(tree_2237)
);
wire [0:0] tree_2238;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2430 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_182),
 .b(tree_87),
 .c(tree_2238)
);
wire [0:0] tree_2239;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2431 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_153),
 .b(tree_331),
 .c(tree_2239)
);
wire [0:0] tree_2240;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2432 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_367),
 .b(tree_54),
 .c(tree_2240)
);
wire [0:0] tree_2241;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2433 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_359),
 .b(tree_12),
 .c(tree_2241)
);
wire [0:0] tree_2242;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2434 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_621),
 .b(1'h0),
 .c(tree_2242)
);
wire [0:0] tree_2243;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2435 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2235),
 .b(tree_2236),
 .c(tree_2243)
);
wire [0:0] tree_2244;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2436 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2237),
 .b(tree_2238),
 .c(tree_2244)
);
wire [0:0] tree_2245;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2437 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2239),
 .b(tree_2240),
 .c(tree_2245)
);
wire [0:0] tree_2246;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2438 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2241),
 .b(tree_2242),
 .c(tree_2246)
);
wire [0:0] tree_2247;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2439 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_700),
 .b(tree_541),
 .c(tree_2247)
);
wire [0:0] tree_2248;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2440 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_459),
 .b(tree_584),
 .c(tree_2248)
);
wire [0:0] tree_2249;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2441 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2243),
 .b(tree_2244),
 .c(tree_2249)
);
wire [0:0] tree_2250;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2442 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2245),
 .b(tree_2246),
 .c(tree_2250)
);
wire [0:0] tree_2251;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2443 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2248),
 .b(tree_2247),
 .c(tree_2251)
);
wire [0:0] tree_2252;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2444 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1234),
 .b(tree_539),
 .c(tree_2252)
);
wire [0:0] tree_2253;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2445 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1203),
 .b(tree_1235),
 .c(tree_2253)
);
wire [0:0] tree_2254;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2446 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_996),
 .b(tree_813),
 .c(tree_2254)
);
wire [0:0] tree_2255;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2447 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2249),
 .b(tree_2250),
 .c(tree_2255)
);
wire [0:0] tree_2256;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2448 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2251),
 .b(tree_2252),
 .c(tree_2256)
);
wire [0:0] tree_2257;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2449 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2253),
 .b(tree_2254),
 .c(tree_2257)
);
wire [0:0] tree_2258;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2450 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2255),
 .b(tree_2256),
 .c(tree_2258)
);
wire [0:0] tree_2259;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2451 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2257),
 .b(1'h0),
 .c(tree_2259)
);
wire [0:0] tree_2260;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2452 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2258),
 .b(tree_2259),
 .c(tree_2260)
);
wire [0:0] tree_2261;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2453 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[7]),
 .b(in[94]),
 .c(tree_2261)
);
wire [0:0] tree_2262;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2454 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[101]),
 .b(in[112]),
 .c(tree_2262)
);
wire [0:0] tree_2263;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2455 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[188]),
 .b(1'h0),
 .c(tree_2263)
);
wire [0:0] tree_2264;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2456 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2262),
 .b(tree_2261),
 .c(tree_2264)
);
wire [0:0] tree_2265;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2457 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2263),
 .b(tree_85),
 .c(tree_2265)
);
wire [0:0] tree_2266;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2458 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_151),
 .b(tree_71),
 .c(tree_2266)
);
wire [0:0] tree_2267;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2459 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_182),
 .b(tree_234),
 .c(tree_2267)
);
wire [0:0] tree_2268;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2460 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_124),
 .b(tree_378),
 .c(tree_2268)
);
wire [0:0] tree_2269;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2461 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_129),
 .b(tree_593),
 .c(tree_2269)
);
wire [0:0] tree_2270;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2462 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_547),
 .b(1'h0),
 .c(tree_2270)
);
wire [0:0] tree_2271;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2463 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2264),
 .b(tree_2265),
 .c(tree_2271)
);
wire [0:0] tree_2272;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2464 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2267),
 .b(tree_2266),
 .c(tree_2272)
);
wire [0:0] tree_2273;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2465 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2268),
 .b(tree_2269),
 .c(tree_2273)
);
wire [0:0] tree_2274;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2466 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2270),
 .b(tree_713),
 .c(tree_2274)
);
wire [0:0] tree_2275;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2467 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_736),
 .b(tree_703),
 .c(tree_2275)
);
wire [0:0] tree_2276;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2468 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_947),
 .b(tree_667),
 .c(tree_2276)
);
wire [0:0] tree_2277;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2469 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_668),
 .b(1'h0),
 .c(tree_2277)
);
wire [0:0] tree_2278;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2470 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2271),
 .b(tree_2272),
 .c(tree_2278)
);
wire [0:0] tree_2279;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2471 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2273),
 .b(tree_2274),
 .c(tree_2279)
);
wire [0:0] tree_2280;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2472 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2275),
 .b(tree_2276),
 .c(tree_2280)
);
wire [0:0] tree_2281;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2473 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1027),
 .b(tree_2277),
 .c(tree_2281)
);
wire [0:0] tree_2282;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2474 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1003),
 .b(tree_643),
 .c(tree_2282)
);
wire [0:0] tree_2283;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2475 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2278),
 .b(tree_2279),
 .c(tree_2283)
);
wire [0:0] tree_2284;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2476 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2280),
 .b(tree_2281),
 .c(tree_2284)
);
wire [0:0] tree_2285;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2477 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2282),
 .b(tree_1855),
 .c(tree_2285)
);
wire [0:0] tree_2286;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2478 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2283),
 .b(tree_2284),
 .c(tree_2286)
);
wire [0:0] tree_2287;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2479 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2285),
 .b(1'h0),
 .c(tree_2287)
);
wire [0:0] tree_2288;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2480 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2286),
 .b(tree_2287),
 .c(tree_2288)
);
wire [0:0] tree_2289;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2481 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[66]),
 .b(in[83]),
 .c(tree_2289)
);
wire [0:0] tree_2290;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2482 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[108]),
 .b(in[168]),
 .c(tree_2290)
);
wire [0:0] tree_2291;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2483 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[191]),
 .b(1'h0),
 .c(tree_2291)
);
wire [0:0] tree_2292;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2484 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2290),
 .b(tree_2289),
 .c(tree_2292)
);
wire [0:0] tree_2293;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2485 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2291),
 .b(tree_42),
 .c(tree_2293)
);
wire [0:0] tree_2294;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2486 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_124),
 .b(tree_162),
 .c(tree_2294)
);
wire [0:0] tree_2295;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2487 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_483),
 .b(tree_490),
 .c(tree_2295)
);
wire [0:0] tree_2296;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2488 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_588),
 .b(tree_510),
 .c(tree_2296)
);
wire [0:0] tree_2297;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2489 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_253),
 .b(tree_594),
 .c(tree_2297)
);
wire [0:0] tree_2298;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2490 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_537),
 .b(1'h0),
 .c(tree_2298)
);
wire [0:0] tree_2299;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2491 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2292),
 .b(tree_2293),
 .c(tree_2299)
);
wire [0:0] tree_2300;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2492 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2294),
 .b(tree_2295),
 .c(tree_2300)
);
wire [0:0] tree_2301;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2493 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2296),
 .b(tree_2297),
 .c(tree_2301)
);
wire [0:0] tree_2302;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2494 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_897),
 .b(tree_2298),
 .c(tree_2302)
);
wire [0:0] tree_2303;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2495 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_749),
 .b(tree_633),
 .c(tree_2303)
);
wire [0:0] tree_2304;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2496 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1041),
 .b(tree_969),
 .c(tree_2304)
);
wire [0:0] tree_2305;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2497 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2299),
 .b(tree_2300),
 .c(tree_2305)
);
wire [0:0] tree_2306;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2498 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2301),
 .b(tree_2302),
 .c(tree_2306)
);
wire [0:0] tree_2307;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2499 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2303),
 .b(tree_2304),
 .c(tree_2307)
);
wire [0:0] tree_2308;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2500 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1503),
 .b(tree_1493),
 .c(tree_2308)
);
wire [0:0] tree_2309;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2501 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1270),
 .b(tree_794),
 .c(tree_2309)
);
wire [0:0] tree_2310;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2502 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1202),
 .b(1'h0),
 .c(tree_2310)
);
wire [0:0] tree_2311;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2503 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2305),
 .b(tree_2306),
 .c(tree_2311)
);
wire [0:0] tree_2312;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2504 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2308),
 .b(tree_2307),
 .c(tree_2312)
);
wire [0:0] tree_2313;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2505 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2309),
 .b(tree_2310),
 .c(tree_2313)
);
wire [0:0] tree_2314;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2506 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2311),
 .b(tree_2312),
 .c(tree_2314)
);
wire [0:0] tree_2315;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2507 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2313),
 .b(1'h0),
 .c(tree_2315)
);
wire [0:0] tree_2316;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2508 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2314),
 .b(tree_2315),
 .c(tree_2316)
);
wire [0:0] tree_2317;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2509 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[26]),
 .b(in[10]),
 .c(tree_2317)
);
wire [0:0] tree_2318;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2510 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[51]),
 .b(in[64]),
 .c(tree_2318)
);
wire [0:0] tree_2319;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2511 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[85]),
 .b(in[89]),
 .c(tree_2319)
);
wire [0:0] tree_2320;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2512 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[97]),
 .b(1'h0),
 .c(tree_2320)
);
wire [0:0] tree_2321;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2513 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2317),
 .b(tree_2318),
 .c(tree_2321)
);
wire [0:0] tree_2322;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2514 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2319),
 .b(tree_2320),
 .c(tree_2322)
);
wire [0:0] tree_2323;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2515 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_85),
 .b(tree_299),
 .c(tree_2323)
);
wire [0:0] tree_2324;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2516 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_164),
 .b(tree_62),
 .c(tree_2324)
);
wire [0:0] tree_2325;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2517 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_335),
 .b(tree_310),
 .c(tree_2325)
);
wire [0:0] tree_2326;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2518 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_34),
 .b(tree_159),
 .c(tree_2326)
);
wire [0:0] tree_2327;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2519 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_471),
 .b(tree_83),
 .c(tree_2327)
);
wire [0:0] tree_2328;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2520 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_146),
 .b(tree_678),
 .c(tree_2328)
);
wire [0:0] tree_2329;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2521 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2321),
 .b(tree_2322),
 .c(tree_2329)
);
wire [0:0] tree_2330;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2522 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2323),
 .b(tree_2324),
 .c(tree_2330)
);
wire [0:0] tree_2331;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2523 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2325),
 .b(tree_2326),
 .c(tree_2331)
);
wire [0:0] tree_2332;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2524 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2327),
 .b(tree_2328),
 .c(tree_2332)
);
wire [0:0] tree_2333;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2525 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_940),
 .b(tree_515),
 .c(tree_2333)
);
wire [0:0] tree_2334;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2526 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_929),
 .b(tree_668),
 .c(tree_2334)
);
wire [0:0] tree_2335;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2527 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2329),
 .b(tree_2330),
 .c(tree_2335)
);
wire [0:0] tree_2336;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2528 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2331),
 .b(tree_2332),
 .c(tree_2336)
);
wire [0:0] tree_2337;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2529 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2333),
 .b(tree_2334),
 .c(tree_2337)
);
wire [0:0] tree_2338;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2530 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_675),
 .b(tree_556),
 .c(tree_2338)
);
wire [0:0] tree_2339;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2531 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_925),
 .b(tree_1272),
 .c(tree_2339)
);
wire [0:0] tree_2340;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2532 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2335),
 .b(tree_2336),
 .c(tree_2340)
);
wire [0:0] tree_2341;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2533 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2337),
 .b(tree_2338),
 .c(tree_2341)
);
wire [0:0] tree_2342;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2534 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2339),
 .b(tree_1499),
 .c(tree_2342)
);
wire [0:0] tree_2343;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2535 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2340),
 .b(tree_2341),
 .c(tree_2343)
);
wire [0:0] tree_2344;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2536 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2342),
 .b(1'h0),
 .c(tree_2344)
);
wire [0:0] tree_2345;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2537 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2343),
 .b(tree_2344),
 .c(tree_2345)
);
wire [0:0] tree_2346;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2538 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[8]),
 .b(in[106]),
 .c(tree_2346)
);
wire [0:0] tree_2347;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2539 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[140]),
 .b(1'h0),
 .c(tree_2347)
);
wire [0:0] tree_2348;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2540 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2346),
 .b(tree_2347),
 .c(tree_2348)
);
wire [0:0] tree_2349;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2541 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_10),
 .b(tree_97),
 .c(tree_2349)
);
wire [0:0] tree_2350;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2542 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_44),
 .b(tree_264),
 .c(tree_2350)
);
wire [0:0] tree_2351;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2543 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_397),
 .b(tree_684),
 .c(tree_2351)
);
wire [0:0] tree_2352;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2544 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_634),
 .b(1'h0),
 .c(tree_2352)
);
wire [0:0] tree_2353;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2545 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2348),
 .b(tree_2349),
 .c(tree_2353)
);
wire [0:0] tree_2354;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2546 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2350),
 .b(tree_2351),
 .c(tree_2354)
);
wire [0:0] tree_2355;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2547 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_711),
 .b(tree_2352),
 .c(tree_2355)
);
wire [0:0] tree_2356;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2548 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_692),
 .b(tree_473),
 .c(tree_2356)
);
wire [0:0] tree_2357;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2549 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_899),
 .b(tree_683),
 .c(tree_2357)
);
wire [0:0] tree_2358;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2550 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_672),
 .b(tree_485),
 .c(tree_2358)
);
wire [0:0] tree_2359;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2551 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_865),
 .b(1'h0),
 .c(tree_2359)
);
wire [0:0] tree_2360;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2552 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2353),
 .b(tree_2354),
 .c(tree_2360)
);
wire [0:0] tree_2361;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2553 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2355),
 .b(tree_2356),
 .c(tree_2361)
);
wire [0:0] tree_2362;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2554 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2357),
 .b(tree_2358),
 .c(tree_2362)
);
wire [0:0] tree_2363;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2555 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1299),
 .b(tree_2359),
 .c(tree_2363)
);
wire [0:0] tree_2364;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2556 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_447),
 .b(tree_949),
 .c(tree_2364)
);
wire [0:0] tree_2365;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2557 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2360),
 .b(tree_2361),
 .c(tree_2365)
);
wire [0:0] tree_2366;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2558 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2362),
 .b(tree_2363),
 .c(tree_2366)
);
wire [0:0] tree_2367;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2559 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2364),
 .b(tree_1919),
 .c(tree_2367)
);
wire [0:0] tree_2368;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2560 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1684),
 .b(1'h0),
 .c(tree_2368)
);
wire [0:0] tree_2369;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2561 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2365),
 .b(tree_2366),
 .c(tree_2369)
);
wire [0:0] tree_2370;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2562 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2367),
 .b(tree_2368),
 .c(tree_2370)
);
wire [0:0] tree_2371;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2563 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2369),
 .b(tree_2370),
 .c(tree_2371)
);
wire [0:0] tree_2372;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2564 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[139]),
 .b(in[95]),
 .c(tree_2372)
);
wire [0:0] tree_2373;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2565 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[155]),
 .b(1'h0),
 .c(tree_2373)
);
wire [0:0] tree_2374;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2566 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2372),
 .b(tree_2373),
 .c(tree_2374)
);
wire [0:0] tree_2375;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2567 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_35),
 .b(tree_163),
 .c(tree_2375)
);
wire [0:0] tree_2376;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2568 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_81),
 .b(tree_376),
 .c(tree_2376)
);
wire [0:0] tree_2377;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2569 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_378),
 .b(tree_133),
 .c(tree_2377)
);
wire [0:0] tree_2378;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2570 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_490),
 .b(tree_510),
 .c(tree_2378)
);
wire [0:0] tree_2379;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2571 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_215),
 .b(tree_599),
 .c(tree_2379)
);
wire [0:0] tree_2380;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2572 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_240),
 .b(1'h0),
 .c(tree_2380)
);
wire [0:0] tree_2381;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2573 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2374),
 .b(tree_2375),
 .c(tree_2381)
);
wire [0:0] tree_2382;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2574 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2376),
 .b(tree_2377),
 .c(tree_2382)
);
wire [0:0] tree_2383;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2575 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2378),
 .b(tree_2379),
 .c(tree_2383)
);
wire [0:0] tree_2384;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2576 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_756),
 .b(tree_2380),
 .c(tree_2384)
);
wire [0:0] tree_2385;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2577 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_418),
 .b(tree_681),
 .c(tree_2385)
);
wire [0:0] tree_2386;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2578 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1015),
 .b(tree_638),
 .c(tree_2386)
);
wire [0:0] tree_2387;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2579 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2381),
 .b(tree_2382),
 .c(tree_2387)
);
wire [0:0] tree_2388;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2580 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2383),
 .b(tree_2384),
 .c(tree_2388)
);
wire [0:0] tree_2389;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2581 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2385),
 .b(tree_2386),
 .c(tree_2389)
);
wire [0:0] tree_2390;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2582 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1234),
 .b(tree_1501),
 .c(tree_2390)
);
wire [0:0] tree_2391;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2583 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1017),
 .b(tree_1117),
 .c(tree_2391)
);
wire [0:0] tree_2392;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2584 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1602),
 .b(1'h0),
 .c(tree_2392)
);
wire [0:0] tree_2393;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2585 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2387),
 .b(tree_2388),
 .c(tree_2393)
);
wire [0:0] tree_2394;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2586 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2389),
 .b(tree_2390),
 .c(tree_2394)
);
wire [0:0] tree_2395;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2587 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2391),
 .b(tree_2392),
 .c(tree_2395)
);
wire [0:0] tree_2396;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2588 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2393),
 .b(tree_2394),
 .c(tree_2396)
);
wire [0:0] tree_2397;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2589 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2395),
 .b(1'h0),
 .c(tree_2397)
);
wire [0:0] tree_2398;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2590 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2396),
 .b(tree_2397),
 .c(tree_2398)
);
wire [0:0] tree_2399;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2591 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[50]),
 .b(in[102]),
 .c(tree_2399)
);
wire [0:0] tree_2400;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2592 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[183]),
 .b(1'h0),
 .c(tree_2400)
);
wire [0:0] tree_2401;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2593 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2399),
 .b(tree_2400),
 .c(tree_2401)
);
wire [0:0] tree_2402;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2594 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_201),
 .b(tree_51),
 .c(tree_2402)
);
wire [0:0] tree_2403;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2595 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_279),
 .b(tree_53),
 .c(tree_2403)
);
wire [0:0] tree_2404;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2596 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_183),
 .b(tree_292),
 .c(tree_2404)
);
wire [0:0] tree_2405;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2597 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_404),
 .b(tree_686),
 .c(tree_2405)
);
wire [0:0] tree_2406;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2598 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_687),
 .b(1'h0),
 .c(tree_2406)
);
wire [0:0] tree_2407;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2599 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2402),
 .b(tree_2401),
 .c(tree_2407)
);
wire [0:0] tree_2408;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2600 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2403),
 .b(tree_2404),
 .c(tree_2408)
);
wire [0:0] tree_2409;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2601 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2405),
 .b(tree_2406),
 .c(tree_2409)
);
wire [0:0] tree_2410;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2602 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_325),
 .b(tree_560),
 .c(tree_2410)
);
wire [0:0] tree_2411;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2603 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_852),
 .b(tree_850),
 .c(tree_2411)
);
wire [0:0] tree_2412;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2604 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_562),
 .b(tree_817),
 .c(tree_2412)
);
wire [0:0] tree_2413;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2605 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_658),
 .b(tree_605),
 .c(tree_2413)
);
wire [0:0] tree_2414;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2606 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_618),
 .b(tree_667),
 .c(tree_2414)
);
wire [0:0] tree_2415;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2607 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2407),
 .b(tree_2408),
 .c(tree_2415)
);
wire [0:0] tree_2416;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2608 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2409),
 .b(tree_2410),
 .c(tree_2416)
);
wire [0:0] tree_2417;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2609 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2411),
 .b(tree_2412),
 .c(tree_2417)
);
wire [0:0] tree_2418;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2610 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2414),
 .b(tree_2413),
 .c(tree_2418)
);
wire [0:0] tree_2419;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2611 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1301),
 .b(tree_375),
 .c(tree_2419)
);
wire [0:0] tree_2420;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2612 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1302),
 .b(1'h0),
 .c(tree_2420)
);
wire [0:0] tree_2421;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2613 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2415),
 .b(tree_2416),
 .c(tree_2421)
);
wire [0:0] tree_2422;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2614 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2417),
 .b(tree_2418),
 .c(tree_2422)
);
wire [0:0] tree_2423;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2615 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2419),
 .b(tree_2420),
 .c(tree_2423)
);
wire [0:0] tree_2424;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2616 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1572),
 .b(1'h0),
 .c(tree_2424)
);
wire [0:0] tree_2425;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2617 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2421),
 .b(tree_2422),
 .c(tree_2425)
);
wire [0:0] tree_2426;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2618 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2423),
 .b(tree_2424),
 .c(tree_2426)
);
wire [0:0] tree_2427;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2619 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2425),
 .b(tree_2426),
 .c(tree_2427)
);
wire [0:0] tree_2428;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2620 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[13]),
 .b(in[91]),
 .c(tree_2428)
);
wire [0:0] tree_2429;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2621 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[158]),
 .b(in[160]),
 .c(tree_2429)
);
wire [0:0] tree_2430;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2622 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2428),
 .b(tree_2429),
 .c(tree_2430)
);
wire [0:0] tree_2431;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2623 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_78),
 .b(tree_305),
 .c(tree_2431)
);
wire [0:0] tree_2432;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2624 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_247),
 .b(tree_412),
 .c(tree_2432)
);
wire [0:0] tree_2433;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2625 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_312),
 .b(tree_251),
 .c(tree_2433)
);
wire [0:0] tree_2434;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2626 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_215),
 .b(tree_632),
 .c(tree_2434)
);
wire [0:0] tree_2435;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2627 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_678),
 .b(tree_445),
 .c(tree_2435)
);
wire [0:0] tree_2436;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2628 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_686),
 .b(tree_687),
 .c(tree_2436)
);
wire [0:0] tree_2437;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2629 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2430),
 .b(tree_2431),
 .c(tree_2437)
);
wire [0:0] tree_2438;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2630 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2433),
 .b(tree_2432),
 .c(tree_2438)
);
wire [0:0] tree_2439;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2631 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2435),
 .b(tree_2434),
 .c(tree_2439)
);
wire [0:0] tree_2440;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2632 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_494),
 .b(tree_2436),
 .c(tree_2440)
);
wire [0:0] tree_2441;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2633 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_698),
 .b(tree_452),
 .c(tree_2441)
);
wire [0:0] tree_2442;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2634 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_351),
 .b(tree_442),
 .c(tree_2442)
);
wire [0:0] tree_2443;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2635 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_511),
 .b(tree_590),
 .c(tree_2443)
);
wire [0:0] tree_2444;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2636 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_93),
 .b(tree_660),
 .c(tree_2444)
);
wire [0:0] tree_2445;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2637 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_646),
 .b(1'h0),
 .c(tree_2445)
);
wire [0:0] tree_2446;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2638 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2437),
 .b(tree_2438),
 .c(tree_2446)
);
wire [0:0] tree_2447;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2639 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2439),
 .b(tree_2440),
 .c(tree_2447)
);
wire [0:0] tree_2448;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2640 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2441),
 .b(tree_2442),
 .c(tree_2448)
);
wire [0:0] tree_2449;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2641 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2443),
 .b(tree_2444),
 .c(tree_2449)
);
wire [0:0] tree_2450;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2642 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1447),
 .b(tree_2445),
 .c(tree_2450)
);
wire [0:0] tree_2451;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2643 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1331),
 .b(tree_1115),
 .c(tree_2451)
);
wire [0:0] tree_2452;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2644 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2446),
 .b(tree_2447),
 .c(tree_2452)
);
wire [0:0] tree_2453;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2645 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2448),
 .b(tree_2449),
 .c(tree_2453)
);
wire [0:0] tree_2454;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2646 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2450),
 .b(tree_2451),
 .c(tree_2454)
);
wire [0:0] tree_2455;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2647 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2452),
 .b(tree_2453),
 .c(tree_2455)
);
wire [0:0] tree_2456;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2648 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2454),
 .b(1'h0),
 .c(tree_2456)
);
wire [0:0] tree_2457;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2649 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2455),
 .b(tree_2456),
 .c(tree_2457)
);
wire [0:0] tree_2458;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2650 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[40]),
 .b(in[35]),
 .c(tree_2458)
);
wire [0:0] tree_2459;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2651 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[93]),
 .b(in[144]),
 .c(tree_2459)
);
wire [0:0] tree_2460;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2652 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[177]),
 .b(1'h0),
 .c(tree_2460)
);
wire [0:0] tree_2461;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2653 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2458),
 .b(tree_2459),
 .c(tree_2461)
);
wire [0:0] tree_2462;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2654 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2460),
 .b(tree_0),
 .c(tree_2462)
);
wire [0:0] tree_2463;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2655 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1),
 .b(tree_2),
 .c(tree_2463)
);
wire [0:0] tree_2464;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2656 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_4),
 .b(tree_3),
 .c(tree_2464)
);
wire [0:0] tree_2465;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2657 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_5),
 .b(tree_8),
 .c(tree_2465)
);
wire [0:0] tree_2466;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2658 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_11),
 .b(tree_12),
 .c(tree_2466)
);
wire [0:0] tree_2467;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2659 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_13),
 .b(tree_17),
 .c(tree_2467)
);
wire [0:0] tree_2468;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2660 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_18),
 .b(tree_19),
 .c(tree_2468)
);
wire [0:0] tree_2469;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2661 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_20),
 .b(1'h0),
 .c(tree_2469)
);
wire [0:0] tree_2470;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2662 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2461),
 .b(tree_2462),
 .c(tree_2470)
);
wire [0:0] tree_2471;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2663 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2464),
 .b(tree_2463),
 .c(tree_2471)
);
wire [0:0] tree_2472;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2664 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2465),
 .b(tree_2466),
 .c(tree_2472)
);
wire [0:0] tree_2473;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2665 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2467),
 .b(tree_2468),
 .c(tree_2473)
);
wire [0:0] tree_2474;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2666 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2469),
 .b(tree_692),
 .c(tree_2474)
);
wire [0:0] tree_2475;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2667 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_694),
 .b(tree_696),
 .c(tree_2475)
);
wire [0:0] tree_2476;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2668 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_700),
 .b(tree_698),
 .c(tree_2476)
);
wire [0:0] tree_2477;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2669 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_703),
 .b(tree_701),
 .c(tree_2477)
);
wire [0:0] tree_2478;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2670 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2470),
 .b(tree_2471),
 .c(tree_2478)
);
wire [0:0] tree_2479;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2671 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2472),
 .b(tree_2473),
 .c(tree_2479)
);
wire [0:0] tree_2480;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2672 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2474),
 .b(tree_2475),
 .c(tree_2480)
);
wire [0:0] tree_2481;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2673 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2476),
 .b(tree_2477),
 .c(tree_2481)
);
wire [0:0] tree_2482;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2674 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1447),
 .b(tree_1445),
 .c(tree_2482)
);
wire [0:0] tree_2483;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2675 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1451),
 .b(tree_1449),
 .c(tree_2483)
);
wire [0:0] tree_2484;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2676 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2478),
 .b(tree_2479),
 .c(tree_2484)
);
wire [0:0] tree_2485;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2677 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2480),
 .b(tree_2481),
 .c(tree_2485)
);
wire [0:0] tree_2486;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2678 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2482),
 .b(tree_2483),
 .c(tree_2486)
);
wire [0:0] tree_2487;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2679 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2484),
 .b(tree_2485),
 .c(tree_2487)
);
wire [0:0] tree_2488;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2680 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2486),
 .b(1'h0),
 .c(tree_2488)
);
wire [0:0] tree_2489;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2681 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2487),
 .b(tree_2488),
 .c(tree_2489)
);
wire [0:0] tree_2490;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2682 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[99]),
 .b(in[137]),
 .c(tree_2490)
);
wire [0:0] tree_2491;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2683 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[156]),
 .b(in[138]),
 .c(tree_2491)
);
wire [0:0] tree_2492;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2684 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2490),
 .b(tree_2491),
 .c(tree_2492)
);
wire [0:0] tree_2493;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2685 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_4),
 .b(tree_32),
 .c(tree_2493)
);
wire [0:0] tree_2494;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2686 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_33),
 .b(tree_34),
 .c(tree_2494)
);
wire [0:0] tree_2495;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2687 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_36),
 .b(tree_11),
 .c(tree_2495)
);
wire [0:0] tree_2496;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2688 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_37),
 .b(tree_45),
 .c(tree_2496)
);
wire [0:0] tree_2497;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2689 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2492),
 .b(tree_2493),
 .c(tree_2497)
);
wire [0:0] tree_2498;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2690 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2494),
 .b(tree_2495),
 .c(tree_2498)
);
wire [0:0] tree_2499;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2691 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2496),
 .b(tree_711),
 .c(tree_2499)
);
wire [0:0] tree_2500;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2692 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_713),
 .b(tree_715),
 .c(tree_2500)
);
wire [0:0] tree_2501;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2693 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_716),
 .b(tree_718),
 .c(tree_2501)
);
wire [0:0] tree_2502;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2694 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_720),
 .b(tree_722),
 .c(tree_2502)
);
wire [0:0] tree_2503;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2695 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_726),
 .b(tree_724),
 .c(tree_2503)
);
wire [0:0] tree_2504;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2696 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_727),
 .b(tree_734),
 .c(tree_2504)
);
wire [0:0] tree_2505;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2697 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2497),
 .b(tree_2498),
 .c(tree_2505)
);
wire [0:0] tree_2506;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2698 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2499),
 .b(tree_2500),
 .c(tree_2506)
);
wire [0:0] tree_2507;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2699 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2502),
 .b(tree_2501),
 .c(tree_2507)
);
wire [0:0] tree_2508;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2700 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2503),
 .b(tree_2504),
 .c(tree_2508)
);
wire [0:0] tree_2509;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2701 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1453),
 .b(tree_1455),
 .c(tree_2509)
);
wire [0:0] tree_2510;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2702 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1457),
 .b(1'h0),
 .c(tree_2510)
);
wire [0:0] tree_2511;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2703 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2505),
 .b(tree_2506),
 .c(tree_2511)
);
wire [0:0] tree_2512;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2704 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2507),
 .b(tree_2508),
 .c(tree_2512)
);
wire [0:0] tree_2513;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2705 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2509),
 .b(tree_2510),
 .c(tree_2513)
);
wire [0:0] tree_2514;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2706 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2511),
 .b(tree_2512),
 .c(tree_2514)
);
wire [0:0] tree_2515;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2707 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2513),
 .b(1'h0),
 .c(tree_2515)
);
wire [0:0] tree_2516;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2708 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2514),
 .b(tree_2515),
 .c(tree_2516)
);
wire [0:0] tree_2517;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2709 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_745),
 .b(1'h0),
 .c(tree_2517)
);
wire [0:0] tree_2518;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2710 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1460),
 .b(tree_2517),
 .c(tree_2518)
);
wire [0:0] tree_2519;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2711 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[3]),
 .b(in[6]),
 .c(tree_2519)
);
wire [0:0] tree_2520;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2712 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[11]),
 .b(in[123]),
 .c(tree_2520)
);
wire [0:0] tree_2521;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2713 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[144]),
 .b(in[186]),
 .c(tree_2521)
);
wire [0:0] tree_2522;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2714 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2519),
 .b(tree_2520),
 .c(tree_2522)
);
wire [0:0] tree_2523;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2715 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2521),
 .b(tree_15),
 .c(tree_2523)
);
wire [0:0] tree_2524;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2716 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_79),
 .b(tree_42),
 .c(tree_2524)
);
wire [0:0] tree_2525;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2717 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_80),
 .b(tree_83),
 .c(tree_2525)
);
wire [0:0] tree_2526;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2718 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_90),
 .b(1'h0),
 .c(tree_2526)
);
wire [0:0] tree_2527;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2719 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2523),
 .b(tree_2522),
 .c(tree_2527)
);
wire [0:0] tree_2528;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2720 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2525),
 .b(tree_2524),
 .c(tree_2528)
);
wire [0:0] tree_2529;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2721 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2526),
 .b(tree_753),
 .c(tree_2529)
);
wire [0:0] tree_2530;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2722 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_755),
 .b(tree_743),
 .c(tree_2530)
);
wire [0:0] tree_2531;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2723 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_756),
 .b(tree_758),
 .c(tree_2531)
);
wire [0:0] tree_2532;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2724 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_768),
 .b(tree_760),
 .c(tree_2532)
);
wire [0:0] tree_2533;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2725 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_773),
 .b(tree_93),
 .c(tree_2533)
);
wire [0:0] tree_2534;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2726 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_774),
 .b(tree_775),
 .c(tree_2534)
);
wire [0:0] tree_2535;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2727 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_780),
 .b(1'h0),
 .c(tree_2535)
);
wire [0:0] tree_2536;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2728 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2527),
 .b(tree_2528),
 .c(tree_2536)
);
wire [0:0] tree_2537;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2729 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2529),
 .b(tree_2530),
 .c(tree_2537)
);
wire [0:0] tree_2538;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2730 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2531),
 .b(tree_2532),
 .c(tree_2538)
);
wire [0:0] tree_2539;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2731 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2533),
 .b(tree_2534),
 .c(tree_2539)
);
wire [0:0] tree_2540;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2732 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2535),
 .b(tree_762),
 .c(tree_2540)
);
wire [0:0] tree_2541;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2733 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_771),
 .b(tree_1462),
 .c(tree_2541)
);
wire [0:0] tree_2542;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2734 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1463),
 .b(1'h0),
 .c(tree_2542)
);
wire [0:0] tree_2543;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2735 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2536),
 .b(tree_2537),
 .c(tree_2543)
);
wire [0:0] tree_2544;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2736 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2538),
 .b(tree_2539),
 .c(tree_2544)
);
wire [0:0] tree_2545;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2737 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2541),
 .b(tree_2540),
 .c(tree_2545)
);
wire [0:0] tree_2546;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2738 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2542),
 .b(1'h0),
 .c(tree_2546)
);
wire [0:0] tree_2547;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2739 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2543),
 .b(tree_2544),
 .c(tree_2547)
);
wire [0:0] tree_2548;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2740 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2545),
 .b(tree_2546),
 .c(tree_2548)
);
wire [0:0] tree_2549;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2741 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2547),
 .b(tree_2548),
 .c(tree_2549)
);
wire [0:0] tree_2550;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2742 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[148]),
 .b(in[6]),
 .c(tree_2550)
);
wire [0:0] tree_2551;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2743 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2550),
 .b(tree_30),
 .c(tree_2551)
);
wire [0:0] tree_2552;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2744 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_1),
 .b(tree_44),
 .c(tree_2552)
);
wire [0:0] tree_2553;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2745 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_32),
 .b(tree_122),
 .c(tree_2553)
);
wire [0:0] tree_2554;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2746 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_123),
 .b(tree_124),
 .c(tree_2554)
);
wire [0:0] tree_2555;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2747 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_125),
 .b(tree_134),
 .c(tree_2555)
);
wire [0:0] tree_2556;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2748 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_135),
 .b(1'h0),
 .c(tree_2556)
);
wire [0:0] tree_2557;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2749 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2551),
 .b(tree_2552),
 .c(tree_2557)
);
wire [0:0] tree_2558;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2750 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2553),
 .b(tree_2554),
 .c(tree_2558)
);
wire [0:0] tree_2559;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2751 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2555),
 .b(tree_2556),
 .c(tree_2559)
);
wire [0:0] tree_2560;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2752 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_796),
 .b(tree_128),
 .c(tree_2560)
);
wire [0:0] tree_2561;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2753 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_798),
 .b(tree_131),
 .c(tree_2561)
);
wire [0:0] tree_2562;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2754 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_802),
 .b(tree_800),
 .c(tree_2562)
);
wire [0:0] tree_2563;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2755 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_804),
 .b(tree_806),
 .c(tree_2563)
);
wire [0:0] tree_2564;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2756 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_808),
 .b(tree_807),
 .c(tree_2564)
);
wire [0:0] tree_2565;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2757 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_809),
 .b(tree_143),
 .c(tree_2565)
);
wire [0:0] tree_2566;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2758 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_810),
 .b(1'h0),
 .c(tree_2566)
);
wire [0:0] tree_2567;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2759 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2557),
 .b(tree_2558),
 .c(tree_2567)
);
wire [0:0] tree_2568;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2760 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2559),
 .b(tree_2560),
 .c(tree_2568)
);
wire [0:0] tree_2569;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2761 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2561),
 .b(tree_2562),
 .c(tree_2569)
);
wire [0:0] tree_2570;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2762 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2563),
 .b(tree_2564),
 .c(tree_2570)
);
wire [0:0] tree_2571;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2763 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2565),
 .b(tree_2566),
 .c(tree_2571)
);
wire [0:0] tree_2572;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2764 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1492),
 .b(tree_813),
 .c(tree_2572)
);
wire [0:0] tree_2573;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2765 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2567),
 .b(tree_2568),
 .c(tree_2573)
);
wire [0:0] tree_2574;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2766 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2569),
 .b(tree_2570),
 .c(tree_2574)
);
wire [0:0] tree_2575;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2767 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2571),
 .b(tree_2572),
 .c(tree_2575)
);
wire [0:0] tree_2576;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2768 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2573),
 .b(tree_2574),
 .c(tree_2576)
);
wire [0:0] tree_2577;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2769 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2575),
 .b(1'h0),
 .c(tree_2577)
);
wire [0:0] tree_2578;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2770 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2576),
 .b(tree_2577),
 .c(tree_2578)
);
wire [0:0] tree_2579;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2771 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[54]),
 .b(in[103]),
 .c(tree_2579)
);
wire [0:0] tree_2580;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2772 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[129]),
 .b(in[135]),
 .c(tree_2580)
);
wire [0:0] tree_2581;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2773 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2579),
 .b(tree_2580),
 .c(tree_2581)
);
wire [0:0] tree_2582;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2774 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_151),
 .b(tree_73),
 .c(tree_2582)
);
wire [0:0] tree_2583;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2775 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_43),
 .b(tree_152),
 .c(tree_2583)
);
wire [0:0] tree_2584;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2776 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_153),
 .b(tree_58),
 .c(tree_2584)
);
wire [0:0] tree_2585;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2777 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_155),
 .b(tree_56),
 .c(tree_2585)
);
wire [0:0] tree_2586;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2778 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2582),
 .b(tree_2581),
 .c(tree_2586)
);
wire [0:0] tree_2587;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2779 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2583),
 .b(tree_2584),
 .c(tree_2587)
);
wire [0:0] tree_2588;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2780 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2585),
 .b(tree_154),
 .c(tree_2588)
);
wire [0:0] tree_2589;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2781 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_814),
 .b(tree_815),
 .c(tree_2589)
);
wire [0:0] tree_2590;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2782 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_817),
 .b(tree_818),
 .c(tree_2590)
);
wire [0:0] tree_2591;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2783 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_824),
 .b(tree_823),
 .c(tree_2591)
);
wire [0:0] tree_2592;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2784 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_825),
 .b(1'h0),
 .c(tree_2592)
);
wire [0:0] tree_2593;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2785 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2586),
 .b(tree_2587),
 .c(tree_2593)
);
wire [0:0] tree_2594;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2786 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2588),
 .b(tree_2589),
 .c(tree_2594)
);
wire [0:0] tree_2595;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2787 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2591),
 .b(tree_2590),
 .c(tree_2595)
);
wire [0:0] tree_2596;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2788 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_821),
 .b(tree_2592),
 .c(tree_2596)
);
wire [0:0] tree_2597;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2789 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1493),
 .b(tree_827),
 .c(tree_2597)
);
wire [0:0] tree_2598;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2790 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1496),
 .b(1'h0),
 .c(tree_2598)
);
wire [0:0] tree_2599;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2791 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2593),
 .b(tree_2594),
 .c(tree_2599)
);
wire [0:0] tree_2600;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2792 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2595),
 .b(tree_2596),
 .c(tree_2600)
);
wire [0:0] tree_2601;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2793 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2597),
 .b(tree_2598),
 .c(tree_2601)
);
wire [0:0] tree_2602;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2794 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1499),
 .b(1'h0),
 .c(tree_2602)
);
wire [0:0] tree_2603;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2795 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2599),
 .b(tree_2600),
 .c(tree_2603)
);
wire [0:0] tree_2604;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2796 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2601),
 .b(tree_2602),
 .c(tree_2604)
);
wire [0:0] tree_2605;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2797 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2603),
 .b(tree_2604),
 .c(tree_2605)
);
wire [0:0] tree_2606;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2798 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[2]),
 .b(in[63]),
 .c(tree_2606)
);
wire [0:0] tree_2607;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2799 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[184]),
 .b(1'h0),
 .c(tree_2607)
);
wire [0:0] tree_2608;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2800 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2606),
 .b(tree_2607),
 .c(tree_2608)
);
wire [0:0] tree_2609;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2801 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_46),
 .b(tree_171),
 .c(tree_2609)
);
wire [0:0] tree_2610;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2802 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_157),
 .b(tree_172),
 .c(tree_2610)
);
wire [0:0] tree_2611;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2803 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_136),
 .b(tree_36),
 .c(tree_2611)
);
wire [0:0] tree_2612;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2804 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2608),
 .b(tree_2609),
 .c(tree_2612)
);
wire [0:0] tree_2613;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2805 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2610),
 .b(tree_2611),
 .c(tree_2613)
);
wire [0:0] tree_2614;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2806 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_753),
 .b(tree_749),
 .c(tree_2614)
);
wire [0:0] tree_2615;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2807 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_836),
 .b(tree_175),
 .c(tree_2615)
);
wire [0:0] tree_2616;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2808 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_811),
 .b(tree_176),
 .c(tree_2616)
);
wire [0:0] tree_2617;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2809 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_179),
 .b(tree_842),
 .c(tree_2617)
);
wire [0:0] tree_2618;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2810 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2612),
 .b(tree_2613),
 .c(tree_2618)
);
wire [0:0] tree_2619;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2811 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2614),
 .b(tree_2615),
 .c(tree_2619)
);
wire [0:0] tree_2620;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2812 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2616),
 .b(tree_2617),
 .c(tree_2620)
);
wire [0:0] tree_2621;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2813 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_839),
 .b(tree_841),
 .c(tree_2621)
);
wire [0:0] tree_2622;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2814 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1501),
 .b(tree_1503),
 .c(tree_2622)
);
wire [0:0] tree_2623;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2815 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1505),
 .b(tree_847),
 .c(tree_2623)
);
wire [0:0] tree_2624;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2816 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2618),
 .b(tree_2619),
 .c(tree_2624)
);
wire [0:0] tree_2625;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2817 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2620),
 .b(tree_2621),
 .c(tree_2625)
);
wire [0:0] tree_2626;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2818 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2622),
 .b(tree_2623),
 .c(tree_2626)
);
wire [0:0] tree_2627;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2819 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2624),
 .b(tree_2625),
 .c(tree_2627)
);
wire [0:0] tree_2628;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2820 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2626),
 .b(1'h0),
 .c(tree_2628)
);
wire [0:0] tree_2629;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2821 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2627),
 .b(tree_2628),
 .c(tree_2629)
);
wire [0:0] tree_2630;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2822 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[101]),
 .b(in[47]),
 .c(tree_2630)
);
wire [0:0] tree_2631;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2823 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[164]),
 .b(in[190]),
 .c(tree_2631)
);
wire [0:0] tree_2632;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2824 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2630),
 .b(tree_2631),
 .c(tree_2632)
);
wire [0:0] tree_2633;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2825 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_61),
 .b(tree_166),
 .c(tree_2633)
);
wire [0:0] tree_2634;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2826 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_211),
 .b(tree_184),
 .c(tree_2634)
);
wire [0:0] tree_2635;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2827 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_215),
 .b(tree_168),
 .c(tree_2635)
);
wire [0:0] tree_2636;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2828 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_218),
 .b(tree_112),
 .c(tree_2636)
);
wire [0:0] tree_2637;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2829 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2632),
 .b(tree_2633),
 .c(tree_2637)
);
wire [0:0] tree_2638;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2830 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2635),
 .b(tree_2634),
 .c(tree_2638)
);
wire [0:0] tree_2639;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2831 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2636),
 .b(tree_177),
 .c(tree_2639)
);
wire [0:0] tree_2640;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2832 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_836),
 .b(tree_863),
 .c(tree_2640)
);
wire [0:0] tree_2641;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2833 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_214),
 .b(tree_217),
 .c(tree_2641)
);
wire [0:0] tree_2642;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2834 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_865),
 .b(tree_220),
 .c(tree_2642)
);
wire [0:0] tree_2643;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2835 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_867),
 .b(tree_872),
 .c(tree_2643)
);
wire [0:0] tree_2644;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2836 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_874),
 .b(tree_873),
 .c(tree_2644)
);
wire [0:0] tree_2645;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2837 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2637),
 .b(tree_2638),
 .c(tree_2645)
);
wire [0:0] tree_2646;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2838 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2640),
 .b(tree_2639),
 .c(tree_2646)
);
wire [0:0] tree_2647;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2839 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2642),
 .b(tree_2641),
 .c(tree_2647)
);
wire [0:0] tree_2648;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2840 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2644),
 .b(tree_2643),
 .c(tree_2648)
);
wire [0:0] tree_2649;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2841 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_876),
 .b(tree_870),
 .c(tree_2649)
);
wire [0:0] tree_2650;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2842 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2645),
 .b(tree_2646),
 .c(tree_2650)
);
wire [0:0] tree_2651;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2843 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2647),
 .b(tree_2648),
 .c(tree_2651)
);
wire [0:0] tree_2652;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2844 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2649),
 .b(tree_1539),
 .c(tree_2652)
);
wire [0:0] tree_2653;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2845 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2650),
 .b(tree_2651),
 .c(tree_2653)
);
wire [0:0] tree_2654;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2846 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2652),
 .b(1'h0),
 .c(tree_2654)
);
wire [0:0] tree_2655;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2847 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2653),
 .b(tree_2654),
 .c(tree_2655)
);
wire [0:0] tree_2656;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2848 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[24]),
 .b(in[68]),
 .c(tree_2656)
);
wire [0:0] tree_2657;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2849 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[69]),
 .b(in[105]),
 .c(tree_2657)
);
wire [0:0] tree_2658;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2850 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[106]),
 .b(1'h0),
 .c(tree_2658)
);
wire [0:0] tree_2659;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2851 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2657),
 .b(tree_2656),
 .c(tree_2659)
);
wire [0:0] tree_2660;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2852 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2658),
 .b(tree_158),
 .c(tree_2660)
);
wire [0:0] tree_2661;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2853 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_235),
 .b(tree_59),
 .c(tree_2661)
);
wire [0:0] tree_2662;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2854 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_253),
 .b(tree_251),
 .c(tree_2662)
);
wire [0:0] tree_2663;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2855 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_259),
 .b(tree_258),
 .c(tree_2663)
);
wire [0:0] tree_2664;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2856 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_45),
 .b(tree_269),
 .c(tree_2664)
);
wire [0:0] tree_2665;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2857 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2659),
 .b(tree_2660),
 .c(tree_2665)
);
wire [0:0] tree_2666;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2858 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2661),
 .b(tree_2662),
 .c(tree_2666)
);
wire [0:0] tree_2667;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2859 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2663),
 .b(tree_2664),
 .c(tree_2667)
);
wire [0:0] tree_2668;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2860 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_889),
 .b(tree_116),
 .c(tree_2668)
);
wire [0:0] tree_2669;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2861 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_257),
 .b(tree_255),
 .c(tree_2669)
);
wire [0:0] tree_2670;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2862 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_891),
 .b(tree_262),
 .c(tree_2670)
);
wire [0:0] tree_2671;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2863 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_892),
 .b(tree_893),
 .c(tree_2671)
);
wire [0:0] tree_2672;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2864 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_268),
 .b(tree_747),
 .c(tree_2672)
);
wire [0:0] tree_2673;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2865 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2665),
 .b(tree_2666),
 .c(tree_2673)
);
wire [0:0] tree_2674;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2866 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2667),
 .b(tree_2668),
 .c(tree_2674)
);
wire [0:0] tree_2675;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2867 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2669),
 .b(tree_2670),
 .c(tree_2675)
);
wire [0:0] tree_2676;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2868 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2671),
 .b(tree_2672),
 .c(tree_2676)
);
wire [0:0] tree_2677;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2869 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1496),
 .b(tree_1569),
 .c(tree_2677)
);
wire [0:0] tree_2678;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2870 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_847),
 .b(1'h0),
 .c(tree_2678)
);
wire [0:0] tree_2679;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2871 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2673),
 .b(tree_2674),
 .c(tree_2679)
);
wire [0:0] tree_2680;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2872 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2675),
 .b(tree_2676),
 .c(tree_2680)
);
wire [0:0] tree_2681;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2873 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2677),
 .b(tree_2678),
 .c(tree_2681)
);
wire [0:0] tree_2682;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2874 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2679),
 .b(tree_2680),
 .c(tree_2682)
);
wire [0:0] tree_2683;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2875 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2681),
 .b(1'h0),
 .c(tree_2683)
);
wire [0:0] tree_2684;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2876 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2682),
 .b(tree_2683),
 .c(tree_2684)
);
wire [0:0] tree_2685;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2877 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[97]),
 .b(in[46]),
 .c(tree_2685)
);
wire [0:0] tree_2686;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2878 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[128]),
 .b(1'h0),
 .c(tree_2686)
);
wire [0:0] tree_2687;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2879 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2685),
 .b(tree_2686),
 .c(tree_2687)
);
wire [0:0] tree_2688;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2880 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_108),
 .b(tree_211),
 .c(tree_2688)
);
wire [0:0] tree_2689;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2881 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_21),
 .b(tree_120),
 .c(tree_2689)
);
wire [0:0] tree_2690;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2882 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_271),
 .b(1'h0),
 .c(tree_2690)
);
wire [0:0] tree_2691;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2883 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2687),
 .b(tree_2688),
 .c(tree_2691)
);
wire [0:0] tree_2692;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2884 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2689),
 .b(tree_2690),
 .c(tree_2692)
);
wire [0:0] tree_2693;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2885 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_897),
 .b(tree_273),
 .c(tree_2693)
);
wire [0:0] tree_2694;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2886 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_262),
 .b(tree_899),
 .c(tree_2694)
);
wire [0:0] tree_2695;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2887 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_907),
 .b(tree_806),
 .c(tree_2695)
);
wire [0:0] tree_2696;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2888 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_727),
 .b(tree_276),
 .c(tree_2696)
);
wire [0:0] tree_2697;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2889 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_909),
 .b(tree_908),
 .c(tree_2697)
);
wire [0:0] tree_2698;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2890 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_867),
 .b(1'h0),
 .c(tree_2698)
);
wire [0:0] tree_2699;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2891 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2691),
 .b(tree_2692),
 .c(tree_2699)
);
wire [0:0] tree_2700;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2892 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2693),
 .b(tree_2694),
 .c(tree_2700)
);
wire [0:0] tree_2701;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2893 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2695),
 .b(tree_2696),
 .c(tree_2701)
);
wire [0:0] tree_2702;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2894 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2697),
 .b(tree_2698),
 .c(tree_2702)
);
wire [0:0] tree_2703;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2895 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_902),
 .b(tree_905),
 .c(tree_2703)
);
wire [0:0] tree_2704;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2896 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_911),
 .b(tree_1451),
 .c(tree_2704)
);
wire [0:0] tree_2705;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2897 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1505),
 .b(1'h0),
 .c(tree_2705)
);
wire [0:0] tree_2706;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2898 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2699),
 .b(tree_2700),
 .c(tree_2706)
);
wire [0:0] tree_2707;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2899 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2701),
 .b(tree_2702),
 .c(tree_2707)
);
wire [0:0] tree_2708;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2900 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2703),
 .b(tree_2704),
 .c(tree_2708)
);
wire [0:0] tree_2709;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2901 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2705),
 .b(tree_1572),
 .c(tree_2709)
);
wire [0:0] tree_2710;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2902 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2706),
 .b(tree_2707),
 .c(tree_2710)
);
wire [0:0] tree_2711;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2903 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2708),
 .b(tree_2709),
 .c(tree_2711)
);
wire [0:0] tree_2712;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2904 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2710),
 .b(tree_2711),
 .c(tree_2712)
);
wire [0:0] tree_2713;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2905 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[1]),
 .b(in[114]),
 .c(tree_2713)
);
wire [0:0] tree_2714;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2906 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[116]),
 .b(in[165]),
 .c(tree_2714)
);
wire [0:0] tree_2715;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2907 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[178]),
 .b(1'h0),
 .c(tree_2715)
);
wire [0:0] tree_2716;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2908 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2714),
 .b(tree_2713),
 .c(tree_2716)
);
wire [0:0] tree_2717;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2909 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2715),
 .b(tree_104),
 .c(tree_2717)
);
wire [0:0] tree_2718;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2910 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_117),
 .b(tree_280),
 .c(tree_2718)
);
wire [0:0] tree_2719;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2911 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_265),
 .b(tree_169),
 .c(tree_2719)
);
wire [0:0] tree_2720;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2912 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_292),
 .b(1'h0),
 .c(tree_2720)
);
wire [0:0] tree_2721;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2913 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2716),
 .b(tree_2717),
 .c(tree_2721)
);
wire [0:0] tree_2722;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2914 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2718),
 .b(tree_2719),
 .c(tree_2722)
);
wire [0:0] tree_2723;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2915 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2720),
 .b(tree_915),
 .c(tree_2723)
);
wire [0:0] tree_2724;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2916 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_287),
 .b(tree_289),
 .c(tree_2724)
);
wire [0:0] tree_2725;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2917 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_291),
 .b(tree_294),
 .c(tree_2725)
);
wire [0:0] tree_2726;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2918 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_296),
 .b(tree_298),
 .c(tree_2726)
);
wire [0:0] tree_2727;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2919 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_917),
 .b(tree_301),
 .c(tree_2727)
);
wire [0:0] tree_2728;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2920 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_825),
 .b(tree_921),
 .c(tree_2728)
);
wire [0:0] tree_2729;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2921 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2721),
 .b(tree_2722),
 .c(tree_2729)
);
wire [0:0] tree_2730;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2922 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2723),
 .b(tree_2724),
 .c(tree_2730)
);
wire [0:0] tree_2731;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2923 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2725),
 .b(tree_2726),
 .c(tree_2731)
);
wire [0:0] tree_2732;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2924 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2727),
 .b(tree_2728),
 .c(tree_2732)
);
wire [0:0] tree_2733;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2925 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_920),
 .b(tree_922),
 .c(tree_2733)
);
wire [0:0] tree_2734;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2926 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1463),
 .b(tree_1573),
 .c(tree_2734)
);
wire [0:0] tree_2735;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2927 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_925),
 .b(1'h0),
 .c(tree_2735)
);
wire [0:0] tree_2736;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2928 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2729),
 .b(tree_2730),
 .c(tree_2736)
);
wire [0:0] tree_2737;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2929 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2731),
 .b(tree_2732),
 .c(tree_2737)
);
wire [0:0] tree_2738;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2930 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2733),
 .b(tree_2734),
 .c(tree_2738)
);
wire [0:0] tree_2739;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2931 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2735),
 .b(1'h0),
 .c(tree_2739)
);
wire [0:0] tree_2740;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2932 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2736),
 .b(tree_2737),
 .c(tree_2740)
);
wire [0:0] tree_2741;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2933 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2738),
 .b(tree_2739),
 .c(tree_2741)
);
wire [0:0] tree_2742;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2934 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2740),
 .b(tree_2741),
 .c(tree_2742)
);
wire [0:0] tree_2743;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2935 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[18]),
 .b(in[21]),
 .c(tree_2743)
);
wire [0:0] tree_2744;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2936 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[93]),
 .b(in[94]),
 .c(tree_2744)
);
wire [0:0] tree_2745;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2937 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[153]),
 .b(in[140]),
 .c(tree_2745)
);
wire [0:0] tree_2746;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2938 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2743),
 .b(tree_2744),
 .c(tree_2746)
);
wire [0:0] tree_2747;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2939 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2745),
 .b(tree_137),
 .c(tree_2747)
);
wire [0:0] tree_2748;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2940 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_275),
 .b(tree_323),
 .c(tree_2748)
);
wire [0:0] tree_2749;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2941 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_41),
 .b(tree_192),
 .c(tree_2749)
);
wire [0:0] tree_2750;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2942 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_326),
 .b(1'h0),
 .c(tree_2750)
);
wire [0:0] tree_2751;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2943 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2746),
 .b(tree_2747),
 .c(tree_2751)
);
wire [0:0] tree_2752;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2944 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2749),
 .b(tree_2748),
 .c(tree_2752)
);
wire [0:0] tree_2753;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2945 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2750),
 .b(tree_325),
 .c(tree_2753)
);
wire [0:0] tree_2754;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2946 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_796),
 .b(tree_932),
 .c(tree_2754)
);
wire [0:0] tree_2755;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2947 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_891),
 .b(tree_329),
 .c(tree_2755)
);
wire [0:0] tree_2756;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2948 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_908),
 .b(tree_935),
 .c(tree_2756)
);
wire [0:0] tree_2757;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2949 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_937),
 .b(1'h0),
 .c(tree_2757)
);
wire [0:0] tree_2758;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2950 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2751),
 .b(tree_2752),
 .c(tree_2758)
);
wire [0:0] tree_2759;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2951 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2753),
 .b(tree_2754),
 .c(tree_2759)
);
wire [0:0] tree_2760;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2952 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2755),
 .b(tree_2756),
 .c(tree_2760)
);
wire [0:0] tree_2761;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2953 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_934),
 .b(tree_2757),
 .c(tree_2761)
);
wire [0:0] tree_2762;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2954 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_333),
 .b(tree_1573),
 .c(tree_2762)
);
wire [0:0] tree_2763;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2955 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1461),
 .b(tree_938),
 .c(tree_2763)
);
wire [0:0] tree_2764;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2956 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1602),
 .b(1'h0),
 .c(tree_2764)
);
wire [0:0] tree_2765;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2957 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2758),
 .b(tree_2759),
 .c(tree_2765)
);
wire [0:0] tree_2766;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2958 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2760),
 .b(tree_2761),
 .c(tree_2766)
);
wire [0:0] tree_2767;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2959 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2762),
 .b(tree_2763),
 .c(tree_2767)
);
wire [0:0] tree_2768;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2960 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2764),
 .b(1'h0),
 .c(tree_2768)
);
wire [0:0] tree_2769;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2961 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2765),
 .b(tree_2766),
 .c(tree_2769)
);
wire [0:0] tree_2770;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2962 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2767),
 .b(tree_2768),
 .c(tree_2770)
);
wire [0:0] tree_2771;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2963 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2769),
 .b(tree_2770),
 .c(tree_2771)
);
wire [0:0] tree_2772;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2964 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[54]),
 .b(in[160]),
 .c(tree_2772)
);
wire [0:0] tree_2773;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2965 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[177]),
 .b(1'h0),
 .c(tree_2773)
);
wire [0:0] tree_2774;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2966 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2772),
 .b(tree_2773),
 .c(tree_2774)
);
wire [0:0] tree_2775;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2967 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_26),
 .b(tree_59),
 .c(tree_2775)
);
wire [0:0] tree_2776;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2968 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_72),
 .b(tree_383),
 .c(tree_2776)
);
wire [0:0] tree_2777;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2969 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_279),
 .b(tree_191),
 .c(tree_2777)
);
wire [0:0] tree_2778;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2970 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_387),
 .b(1'h0),
 .c(tree_2778)
);
wire [0:0] tree_2779;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2971 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2774),
 .b(tree_2775),
 .c(tree_2779)
);
wire [0:0] tree_2780;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2972 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2776),
 .b(tree_2777),
 .c(tree_2780)
);
wire [0:0] tree_2781;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2973 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2778),
 .b(tree_743),
 .c(tree_2781)
);
wire [0:0] tree_2782;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2974 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_385),
 .b(tree_370),
 .c(tree_2782)
);
wire [0:0] tree_2783;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2975 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_966),
 .b(tree_389),
 .c(tree_2783)
);
wire [0:0] tree_2784;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2976 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_946),
 .b(tree_391),
 .c(tree_2784)
);
wire [0:0] tree_2785;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2977 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_968),
 .b(tree_276),
 .c(tree_2785)
);
wire [0:0] tree_2786;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2978 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_394),
 .b(tree_969),
 .c(tree_2786)
);
wire [0:0] tree_2787;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2979 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_970),
 .b(1'h0),
 .c(tree_2787)
);
wire [0:0] tree_2788;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2980 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2779),
 .b(tree_2780),
 .c(tree_2788)
);
wire [0:0] tree_2789;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2981 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2781),
 .b(tree_2782),
 .c(tree_2789)
);
wire [0:0] tree_2790;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2982 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2783),
 .b(tree_2784),
 .c(tree_2790)
);
wire [0:0] tree_2791;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2983 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2785),
 .b(tree_2786),
 .c(tree_2791)
);
wire [0:0] tree_2792;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2984 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2787),
 .b(tree_972),
 .c(tree_2792)
);
wire [0:0] tree_2793;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2985 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2788),
 .b(tree_2789),
 .c(tree_2793)
);
wire [0:0] tree_2794;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2986 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2790),
 .b(tree_2791),
 .c(tree_2794)
);
wire [0:0] tree_2795;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2987 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2792),
 .b(tree_1684),
 .c(tree_2795)
);
wire [0:0] tree_2796;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2988 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2793),
 .b(tree_2794),
 .c(tree_2796)
);
wire [0:0] tree_2797;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2989 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2795),
 .b(1'h0),
 .c(tree_2797)
);
wire [0:0] tree_2798;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2990 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2796),
 .b(tree_2797),
 .c(tree_2798)
);
wire [0:0] tree_2799;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2991 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[43]),
 .b(in[21]),
 .c(tree_2799)
);
wire [0:0] tree_2800;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2992 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[83]),
 .b(in[133]),
 .c(tree_2800)
);
wire [0:0] tree_2801;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2993 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[147]),
 .b(1'h0),
 .c(tree_2801)
);
wire [0:0] tree_2802;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2994 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2799),
 .b(tree_2800),
 .c(tree_2802)
);
wire [0:0] tree_2803;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2995 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_165),
 .b(tree_2801),
 .c(tree_2803)
);
wire [0:0] tree_2804;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_2996 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_163),
 .b(tree_103),
 .c(tree_2804)
);
wire [0:0] tree_2805;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2997 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_299),
 .b(tree_263),
 .c(tree_2805)
);
wire [0:0] tree_2806;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2998 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_72),
 .b(tree_74),
 .c(tree_2806)
);
wire [0:0] tree_2807;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_2999 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_361),
 .b(tree_227),
 .c(tree_2807)
);
wire [0:0] tree_2808;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3000 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_250),
 .b(tree_258),
 .c(tree_2808)
);
wire [0:0] tree_2809;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3001 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_445),
 .b(1'h0),
 .c(tree_2809)
);
wire [0:0] tree_2810;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3002 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2802),
 .b(tree_2803),
 .c(tree_2810)
);
wire [0:0] tree_2811;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3003 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2805),
 .b(tree_2804),
 .c(tree_2811)
);
wire [0:0] tree_2812;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3004 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2806),
 .b(tree_2807),
 .c(tree_2812)
);
wire [0:0] tree_2813;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3005 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2808),
 .b(tree_2809),
 .c(tree_2813)
);
wire [0:0] tree_2814;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3006 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_434),
 .b(tree_436),
 .c(tree_2814)
);
wire [0:0] tree_2815;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3007 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_438),
 .b(tree_440),
 .c(tree_2815)
);
wire [0:0] tree_2816;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3008 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_442),
 .b(tree_852),
 .c(tree_2816)
);
wire [0:0] tree_2817;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3009 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_444),
 .b(tree_179),
 .c(tree_2817)
);
wire [0:0] tree_2818;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3010 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2810),
 .b(tree_2811),
 .c(tree_2818)
);
wire [0:0] tree_2819;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3011 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2812),
 .b(tree_2813),
 .c(tree_2819)
);
wire [0:0] tree_2820;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3012 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2814),
 .b(tree_2815),
 .c(tree_2820)
);
wire [0:0] tree_2821;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3013 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2817),
 .b(tree_2816),
 .c(tree_2821)
);
wire [0:0] tree_2822;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3014 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_989),
 .b(tree_986),
 .c(tree_2822)
);
wire [0:0] tree_2823;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3015 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_447),
 .b(tree_860),
 .c(tree_2823)
);
wire [0:0] tree_2824;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3016 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_333),
 .b(tree_1742),
 .c(tree_2824)
);
wire [0:0] tree_2825;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3017 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2818),
 .b(tree_2819),
 .c(tree_2825)
);
wire [0:0] tree_2826;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3018 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2820),
 .b(tree_2821),
 .c(tree_2826)
);
wire [0:0] tree_2827;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3019 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2822),
 .b(tree_2823),
 .c(tree_2827)
);
wire [0:0] tree_2828;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3020 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2824),
 .b(1'h0),
 .c(tree_2828)
);
wire [0:0] tree_2829;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3021 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2825),
 .b(tree_2826),
 .c(tree_2829)
);
wire [0:0] tree_2830;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3022 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2827),
 .b(tree_2828),
 .c(tree_2830)
);
wire [0:0] tree_2831;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3023 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2829),
 .b(tree_2830),
 .c(tree_2831)
);
wire [0:0] tree_2832;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3024 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[111]),
 .b(in[25]),
 .c(tree_2832)
);
wire [0:0] tree_2833;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3025 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[183]),
 .b(1'h0),
 .c(tree_2833)
);
wire [0:0] tree_2834;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3026 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2832),
 .b(tree_2833),
 .c(tree_2834)
);
wire [0:0] tree_2835;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3027 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_167),
 .b(tree_462),
 .c(tree_2835)
);
wire [0:0] tree_2836;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3028 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_342),
 .b(tree_510),
 .c(tree_2836)
);
wire [0:0] tree_2837;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3029 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_135),
 .b(tree_236),
 .c(tree_2837)
);
wire [0:0] tree_2838;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3030 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2834),
 .b(tree_2835),
 .c(tree_2838)
);
wire [0:0] tree_2839;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3031 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2836),
 .b(tree_2837),
 .c(tree_2839)
);
wire [0:0] tree_2840;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3032 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_766),
 .b(tree_511),
 .c(tree_2840)
);
wire [0:0] tree_2841;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3033 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_469),
 .b(tree_818),
 .c(tree_2841)
);
wire [0:0] tree_2842;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3034 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_513),
 .b(tree_298),
 .c(tree_2842)
);
wire [0:0] tree_2843;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3035 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_509),
 .b(1'h0),
 .c(tree_2843)
);
wire [0:0] tree_2844;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3036 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2838),
 .b(tree_2839),
 .c(tree_2844)
);
wire [0:0] tree_2845;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3037 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2841),
 .b(tree_2840),
 .c(tree_2845)
);
wire [0:0] tree_2846;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3038 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2843),
 .b(tree_2842),
 .c(tree_2846)
);
wire [0:0] tree_2847;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3039 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_983),
 .b(tree_1455),
 .c(tree_2847)
);
wire [0:0] tree_2848;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3040 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2844),
 .b(tree_2845),
 .c(tree_2848)
);
wire [0:0] tree_2849;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3041 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2846),
 .b(tree_2847),
 .c(tree_2849)
);
wire [0:0] tree_2850;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3042 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1853),
 .b(tree_1855),
 .c(tree_2850)
);
wire [0:0] tree_2851;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3043 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1539),
 .b(1'h0),
 .c(tree_2851)
);
wire [0:0] tree_2852;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3044 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2848),
 .b(tree_2849),
 .c(tree_2852)
);
wire [0:0] tree_2853;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3045 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2850),
 .b(tree_2851),
 .c(tree_2853)
);
wire [0:0] tree_2854;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3046 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2852),
 .b(tree_2853),
 .c(tree_2854)
);
wire [0:0] tree_2855;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3047 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[39]),
 .b(in[60]),
 .c(tree_2855)
);
wire [0:0] tree_2856;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3048 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[123]),
 .b(1'h0),
 .c(tree_2856)
);
wire [0:0] tree_2857;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3049 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2855),
 .b(tree_2856),
 .c(tree_2857)
);
wire [0:0] tree_2858;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3050 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_166),
 .b(tree_138),
 .c(tree_2858)
);
wire [0:0] tree_2859;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3051 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_544),
 .b(tree_8),
 .c(tree_2859)
);
wire [0:0] tree_2860;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3052 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_367),
 .b(tree_547),
 .c(tree_2860)
);
wire [0:0] tree_2861;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3053 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_550),
 .b(tree_409),
 .c(tree_2861)
);
wire [0:0] tree_2862;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3054 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_75),
 .b(1'h0),
 .c(tree_2862)
);
wire [0:0] tree_2863;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3055 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2857),
 .b(tree_2858),
 .c(tree_2863)
);
wire [0:0] tree_2864;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3056 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2859),
 .b(tree_2860),
 .c(tree_2864)
);
wire [0:0] tree_2865;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3057 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2861),
 .b(tree_2862),
 .c(tree_2865)
);
wire [0:0] tree_2866;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3058 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_753),
 .b(tree_425),
 .c(tree_2866)
);
wire [0:0] tree_2867;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3059 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_546),
 .b(tree_438),
 .c(tree_2867)
);
wire [0:0] tree_2868;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3060 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_814),
 .b(tree_294),
 .c(tree_2868)
);
wire [0:0] tree_2869;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3061 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_552),
 .b(tree_549),
 .c(tree_2869)
);
wire [0:0] tree_2870;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3062 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_478),
 .b(tree_554),
 .c(tree_2870)
);
wire [0:0] tree_2871;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3063 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1031),
 .b(1'h0),
 .c(tree_2871)
);
wire [0:0] tree_2872;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3064 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2863),
 .b(tree_2864),
 .c(tree_2872)
);
wire [0:0] tree_2873;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3065 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2865),
 .b(tree_2866),
 .c(tree_2873)
);
wire [0:0] tree_2874;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3066 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2867),
 .b(tree_2868),
 .c(tree_2874)
);
wire [0:0] tree_2875;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3067 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2869),
 .b(tree_2870),
 .c(tree_2875)
);
wire [0:0] tree_2876;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3068 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_986),
 .b(tree_2871),
 .c(tree_2876)
);
wire [0:0] tree_2877;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3069 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1030),
 .b(tree_556),
 .c(tree_2877)
);
wire [0:0] tree_2878;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3070 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2872),
 .b(tree_2873),
 .c(tree_2878)
);
wire [0:0] tree_2879;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3071 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2874),
 .b(tree_2875),
 .c(tree_2879)
);
wire [0:0] tree_2880;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3072 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2876),
 .b(tree_2877),
 .c(tree_2880)
);
wire [0:0] tree_2881;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3073 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_1919),
 .b(1'h0),
 .c(tree_2881)
);
wire [0:0] tree_2882;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3074 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2878),
 .b(tree_2879),
 .c(tree_2882)
);
wire [0:0] tree_2883;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3075 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2880),
 .b(tree_2881),
 .c(tree_2883)
);
wire [0:0] tree_2884;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3076 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2882),
 .b(tree_2883),
 .c(tree_2884)
);
wire [0:0] tree_2885;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3077 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[91]),
 .b(1'h0),
 .c(tree_2885)
);
wire [0:0] tree_2886;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3078 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2885),
 .b(tree_96),
 .c(tree_2886)
);
wire [0:0] tree_2887;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3079 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_274),
 .b(tree_26),
 .c(tree_2887)
);
wire [0:0] tree_2888;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3080 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_153),
 .b(tree_69),
 .c(tree_2888)
);
wire [0:0] tree_2889;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3081 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_577),
 .b(tree_125),
 .c(tree_2889)
);
wire [0:0] tree_2890;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3082 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_322),
 .b(tree_579),
 .c(tree_2890)
);
wire [0:0] tree_2891;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3083 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_210),
 .b(tree_580),
 .c(tree_2891)
);
wire [0:0] tree_2892;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3084 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_90),
 .b(tree_523),
 .c(tree_2892)
);
wire [0:0] tree_2893;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3085 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2887),
 .b(tree_2886),
 .c(tree_2893)
);
wire [0:0] tree_2894;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3086 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2889),
 .b(tree_2888),
 .c(tree_2894)
);
wire [0:0] tree_2895;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3087 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2890),
 .b(tree_2891),
 .c(tree_2895)
);
wire [0:0] tree_2896;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3088 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2892),
 .b(tree_576),
 .c(tree_2896)
);
wire [0:0] tree_2897;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3089 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_438),
 .b(tree_291),
 .c(tree_2897)
);
wire [0:0] tree_2898;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3090 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_578),
 .b(tree_255),
 .c(tree_2898)
);
wire [0:0] tree_2899;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3091 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_582),
 .b(tree_346),
 .c(tree_2899)
);
wire [0:0] tree_2900;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3092 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_1036),
 .b(tree_480),
 .c(tree_2900)
);
wire [0:0] tree_2901;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3093 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_888),
 .b(1'h0),
 .c(tree_2901)
);
wire [0:0] tree_2902;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3094 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2893),
 .b(tree_2894),
 .c(tree_2902)
);
wire [0:0] tree_2903;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3095 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2895),
 .b(tree_2896),
 .c(tree_2903)
);
wire [0:0] tree_2904;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3096 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2897),
 .b(tree_2898),
 .c(tree_2904)
);
wire [0:0] tree_2905;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3097 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2899),
 .b(tree_2900),
 .c(tree_2905)
);
wire [0:0] tree_2906;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3098 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2901),
 .b(tree_1018),
 .c(tree_2906)
);
wire [0:0] tree_2907;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3099 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2902),
 .b(tree_2903),
 .c(tree_2907)
);
wire [0:0] tree_2908;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3100 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2904),
 .b(tree_2905),
 .c(tree_2908)
);
wire [0:0] tree_2909;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3101 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2906),
 .b(tree_2518),
 .c(tree_2909)
);
wire [0:0] tree_2910;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3102 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2907),
 .b(tree_2908),
 .c(tree_2910)
);
wire [0:0] tree_2911;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3103 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2909),
 .b(1'h0),
 .c(tree_2911)
);
wire [0:0] tree_2912;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3104 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2910),
 .b(tree_2911),
 .c(tree_2912)
);
wire [0:0] tree_2913;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3105 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[58]),
 .b(in[76]),
 .c(tree_2913)
);
wire [0:0] tree_2914;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3106 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[104]),
 .b(in[152]),
 .c(tree_2914)
);
wire [0:0] tree_2915;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3107 (
 .clk(clock),
 .reset(resets[0]),
 .a(in[158]),
 .b(1'h0),
 .c(tree_2915)
);
wire [0:0] tree_2916;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3108 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_2913),
 .b(tree_2914),
 .c(tree_2916)
);
wire [0:0] tree_2917;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3109 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_6),
 .b(tree_2915),
 .c(tree_2917)
);
wire [0:0] tree_2918;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3110 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_21),
 .b(tree_58),
 .c(tree_2918)
);
wire [0:0] tree_2919;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3111 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_60),
 .b(tree_63),
 .c(tree_2919)
);
wire [0:0] tree_2920;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3112 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_65),
 .b(tree_66),
 .c(tree_2920)
);
wire [0:0] tree_2921;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3113 (
 .clk(clock),
 .reset(resets[1]),
 .a(tree_75),
 .b(tree_67),
 .c(tree_2921)
);
wire [0:0] tree_2922;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3114 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2917),
 .b(tree_2916),
 .c(tree_2922)
);
wire [0:0] tree_2923;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3115 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2918),
 .b(tree_2919),
 .c(tree_2923)
);
wire [0:0] tree_2924;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3116 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_2920),
 .b(tree_2921),
 .c(tree_2924)
);
wire [0:0] tree_2925;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3117 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_735),
 .b(tree_700),
 .c(tree_2925)
);
wire [0:0] tree_2926;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3118 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_738),
 .b(tree_736),
 .c(tree_2926)
);
wire [0:0] tree_2927;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3119 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_740),
 .b(tree_739),
 .c(tree_2927)
);
wire [0:0] tree_2928;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3120 (
 .clk(clock),
 .reset(resets[2]),
 .a(tree_741),
 .b(tree_747),
 .c(tree_2928)
);
wire [0:0] tree_2929;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3121 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2922),
 .b(tree_2923),
 .c(tree_2929)
);
wire [0:0] tree_2930;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3122 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2924),
 .b(tree_2925),
 .c(tree_2930)
);
wire [0:0] tree_2931;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3123 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2926),
 .b(tree_2927),
 .c(tree_2931)
);
wire [0:0] tree_2932;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3124 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_2928),
 .b(tree_1445),
 .c(tree_2932)
);
wire [0:0] tree_2933;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3125 (
 .clk(clock),
 .reset(resets[3]),
 .a(tree_1461),
 .b(1'h0),
 .c(tree_2933)
);
wire [0:0] tree_2934;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3126 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2929),
 .b(tree_2930),
 .c(tree_2934)
);
wire [0:0] tree_2935;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3127 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2931),
 .b(tree_2932),
 .c(tree_2935)
);
wire [0:0] tree_2936;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3128 (
 .clk(clock),
 .reset(resets[4]),
 .a(tree_2933),
 .b(tree_2518),
 .c(tree_2936)
);
wire [0:0] tree_2937;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3129 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2934),
 .b(tree_2935),
 .c(tree_2937)
);
wire [0:0] tree_2938;
serial_adder #(
  .neg_b(1),
  .BW(1)
) op_3130 (
 .clk(clock),
 .reset(resets[5]),
 .a(tree_2936),
 .b(1'h0),
 .c(tree_2938)
);
wire [0:0] tree_2939;
serial_adder #(
  .neg_b(0),
  .BW(1)
) op_3131 (
 .clk(clock),
 .reset(resets[6]),
 .a(tree_2937),
 .b(tree_2938),
 .c(tree_2939)
);
assign out[0] = tree_2489;
assign out[1] = tree_2516;
assign out[2] = tree_2939;
assign out[3] = tree_2549;
assign out[4] = tree_1490;
assign out[5] = tree_2578;
assign out[6] = tree_2605;
assign out[7] = tree_2629;
assign out[8] = tree_1537;
assign out[9] = tree_2655;
assign out[10] = tree_1567;
assign out[11] = tree_2684;
assign out[12] = tree_2712;
assign out[13] = tree_2742;
assign out[14] = tree_1601;
assign out[15] = tree_2771;
assign out[16] = tree_1625;
assign out[17] = tree_1654;
assign out[18] = tree_1682;
assign out[19] = tree_2798;
assign out[20] = tree_1713;
assign out[21] = tree_1741;
assign out[22] = tree_2831;
assign out[23] = tree_1767;
assign out[24] = tree_1794;
assign out[25] = tree_1823;
assign out[26] = tree_1850;
assign out[27] = tree_2854;
assign out[28] = tree_1885;
assign out[29] = tree_1916;
assign out[30] = tree_2884;
assign out[31] = tree_1948;
assign out[32] = tree_1972;
assign out[33] = tree_2912;
assign out[34] = tree_1999;
assign out[35] = tree_2030;
assign out[36] = tree_2059;
assign out[37] = tree_2088;
assign out[38] = tree_1072;
assign out[39] = tree_1103;
assign out[40] = tree_2117;
assign out[41] = tree_2145;
assign out[42] = tree_2174;
assign out[43] = tree_1145;
assign out[44] = tree_1172;
assign out[45] = tree_1199;
assign out[46] = tree_2199;
assign out[47] = tree_2230;
assign out[48] = tree_1231;
assign out[49] = tree_2260;
assign out[50] = tree_2288;
assign out[51] = tree_1268;
assign out[52] = tree_2316;
assign out[53] = tree_2345;
assign out[54] = tree_1297;
assign out[55] = tree_2371;
assign out[56] = tree_2398;
assign out[57] = tree_2427;
assign out[58] = tree_1330;
assign out[59] = tree_2457;
assign out[60] = tree_1360;
assign out[61] = tree_1388;
assign out[62] = tree_1418;
assign out[63] = tree_1443;
always @( posedge clock ) begin

end
endmodule
