localparam D3_IN_SIZE = 1;
localparam D3_BW_W = 16;
localparam D3_SHIFT = 6;
localparam LOG2_D3_CYC = 7;
localparam D3_CYC = 128;
localparam D3_CH = 4;
reg [LOG2_D3_CYC-1:0] d3_cntr;
wire [D3_CH-1:0][D3_IN_SIZE*D3_BW_W-1:0] dw_3;
reg [D3_CYC-1:0][D3_IN_SIZE*D3_BW_W-1:0] dw_3_0 = { 16'hfff1, 16'h000b, 16'hfffb, 16'hfff9, 16'h0000, 16'h0003, 16'hfffa, 16'hfff3, 16'hfff8, 16'hfff2, 16'hfff2, 16'h0008, 16'h0006, 16'h0006, 16'hfff7, 16'h0007, 16'hfff8, 16'h0002, 16'hfff5, 16'h0010, 16'h0009, 16'hfff6, 16'hfff2, 16'h000d, 16'h000a, 16'hfffe, 16'hffff, 16'h000b, 16'h0004, 16'hfff7, 16'h0012, 16'h0002, 16'h000d, 16'hfffb, 16'hfff6, 16'h0004, 16'hfff5, 16'h000f, 16'hfff2, 16'hffff, 16'h0007, 16'h000d, 16'h0000, 16'h0000, 16'hfff3, 16'h000e, 16'h0009, 16'hfffc, 16'hfff2, 16'h0008, 16'h000e, 16'h0006, 16'h0009, 16'hffed, 16'hfff1, 16'hfffc, 16'hfff6, 16'h0005, 16'hfff1, 16'hfffb, 16'hfffe, 16'hfffb, 16'h0009, 16'hfff0, 16'hfff3, 16'hfff7, 16'hfff4, 16'hfffc, 16'hffff, 16'hfff3, 16'hfff9, 16'hffff, 16'hfffe, 16'hfff2, 16'hfffd, 16'hfff5, 16'hfff6, 16'hfff1, 16'h0003, 16'hfffd, 16'h000c, 16'h0003, 16'h0000, 16'hfffa, 16'h0012, 16'hfff0, 16'h0001, 16'hfffa, 16'h0006, 16'hfff9, 16'h0012, 16'hfffe, 16'hfffd, 16'h000f, 16'h0005, 16'h0011, 16'hfff5, 16'h0000, 16'h0004, 16'hfff1, 16'h0010, 16'hfff2, 16'h0008, 16'hffef, 16'h0003, 16'h000f, 16'hfff1, 16'h0010, 16'h0001, 16'h0005, 16'hfffd, 16'hfffb, 16'hfffd, 16'hfff7, 16'hfff7, 16'h000e, 16'h0008, 16'h0006, 16'hfff7, 16'h000c, 16'h000e, 16'h000b, 16'h0015, 16'h0004, 16'h0000, 16'hfffb, 16'hfff0, 16'hfffa };
assign dw_3[0] = dw_3_0[d3_cntr];
reg [D3_CYC-1:0][D3_IN_SIZE*D3_BW_W-1:0] dw_3_1 = { 16'h000b, 16'h0007, 16'h000b, 16'hfff8, 16'h0001, 16'hfff5, 16'h0007, 16'h000c, 16'h0012, 16'hfffc, 16'h000c, 16'hfff2, 16'h0002, 16'h000d, 16'hfffc, 16'h0000, 16'h000b, 16'h0004, 16'hfff6, 16'h000b, 16'h0010, 16'h000e, 16'hfffd, 16'h0002, 16'h0011, 16'hfff6, 16'h0002, 16'hfffa, 16'h0000, 16'hfffb, 16'hfffd, 16'hfff7, 16'hfffc, 16'h000d, 16'h000b, 16'h000e, 16'hfff1, 16'hfff5, 16'h0009, 16'h0007, 16'hfffc, 16'h0006, 16'hfffd, 16'h000b, 16'hfff3, 16'hfff0, 16'h0008, 16'hfff3, 16'h0012, 16'hfffc, 16'hfff7, 16'hfff8, 16'hfff5, 16'h000e, 16'hfffd, 16'hfffd, 16'hfff3, 16'hfff5, 16'hfff5, 16'hfff8, 16'h0005, 16'hfff4, 16'hfffd, 16'hfff9, 16'hfff5, 16'hfff1, 16'h000b, 16'hfff1, 16'h0008, 16'h000e, 16'h0005, 16'h0007, 16'h000c, 16'h000d, 16'h000f, 16'h0007, 16'hfffd, 16'h0002, 16'hfffd, 16'hfff3, 16'hfff5, 16'h0003, 16'hffff, 16'hffef, 16'hfffa, 16'h000d, 16'hfffb, 16'h0001, 16'hfffe, 16'h0003, 16'h0003, 16'h0004, 16'h000d, 16'h0008, 16'hfff8, 16'hffef, 16'hfff3, 16'hfffd, 16'hfff3, 16'hfff2, 16'hfffc, 16'hfff7, 16'hfffc, 16'h0001, 16'h0012, 16'h0001, 16'h0002, 16'h000c, 16'hffff, 16'h0004, 16'hffff, 16'h000d, 16'h0010, 16'h0007, 16'h0003, 16'h0000, 16'h000e, 16'hfff3, 16'h0005, 16'hfff8, 16'h0002, 16'hfffc, 16'h0006, 16'h0005, 16'h0000, 16'h000b, 16'h0002, 16'hffef };
assign dw_3[1] = dw_3_1[d3_cntr];
reg [D3_CYC-1:0][D3_IN_SIZE*D3_BW_W-1:0] dw_3_2 = { 16'h0009, 16'hfff2, 16'h0006, 16'h0008, 16'hfff6, 16'h000e, 16'hfff8, 16'h0001, 16'hfffc, 16'hfff4, 16'h0005, 16'hffff, 16'h0001, 16'hffff, 16'h0003, 16'hfffb, 16'hfffb, 16'h000d, 16'h0006, 16'hfff6, 16'h0003, 16'hfff5, 16'h000e, 16'h0003, 16'hfffb, 16'hfffa, 16'h000f, 16'h0008, 16'h000a, 16'hffff, 16'hfff6, 16'hfff7, 16'hfff6, 16'hffef, 16'h0001, 16'hfff6, 16'h000c, 16'h0007, 16'h000c, 16'h0002, 16'hfff2, 16'h000b, 16'h000a, 16'hfff4, 16'h0006, 16'hfff8, 16'hfffd, 16'h000d, 16'h0002, 16'h0002, 16'h0004, 16'h000c, 16'h000a, 16'hfffe, 16'h000a, 16'hfff9, 16'h000f, 16'hfffa, 16'hfff3, 16'h0010, 16'hfffd, 16'h0009, 16'h0002, 16'h0001, 16'h000e, 16'h0011, 16'h0011, 16'h0007, 16'h000a, 16'hfffc, 16'hfffc, 16'h0010, 16'h0003, 16'h0004, 16'hfffc, 16'hfff3, 16'hffff, 16'hfff3, 16'hffff, 16'hfff8, 16'hfff8, 16'h000b, 16'h0008, 16'hfffe, 16'h0006, 16'hffff, 16'h0007, 16'h0008, 16'h000e, 16'hfffc, 16'h0009, 16'hfff2, 16'hfff8, 16'h000a, 16'h0005, 16'hfffc, 16'h000c, 16'hfff7, 16'h0005, 16'h000c, 16'h0004, 16'h0000, 16'hfff9, 16'h000b, 16'h000a, 16'hfffb, 16'hfffe, 16'hfff4, 16'hfff9, 16'hfffd, 16'hffef, 16'h0000, 16'h0008, 16'hfff3, 16'hfffe, 16'hfffc, 16'h0000, 16'hffff, 16'h0009, 16'hfffc, 16'hffec, 16'h0005, 16'h0002, 16'hfffb, 16'hfff5, 16'hfffb, 16'h000d, 16'hfffc };
assign dw_3[2] = dw_3_2[d3_cntr];
reg [D3_CYC-1:0][D3_IN_SIZE*D3_BW_W-1:0] dw_3_3 = { 16'hfff2, 16'hfff2, 16'hfff5, 16'hfff9, 16'hfff3, 16'h0004, 16'hfff7, 16'hfff9, 16'hfffa, 16'h0011, 16'h0008, 16'hfff8, 16'hfffd, 16'hfffb, 16'hfff6, 16'hfff2, 16'h0007, 16'h0007, 16'hfffb, 16'hfffe, 16'h0004, 16'h0006, 16'hfff3, 16'hfffb, 16'h0005, 16'h000b, 16'h000a, 16'hfffa, 16'hfff3, 16'h000e, 16'h000f, 16'h000c, 16'hfff3, 16'h0000, 16'h0008, 16'hfff6, 16'h000c, 16'h0008, 16'hfff7, 16'h000e, 16'hfff8, 16'hfff0, 16'hfff9, 16'h0005, 16'h0009, 16'h0006, 16'h000c, 16'h000b, 16'hfffc, 16'hfff9, 16'h0004, 16'hfffe, 16'hfff4, 16'h0008, 16'hffff, 16'h000d, 16'hfff8, 16'hffff, 16'h0000, 16'hfff7, 16'h000a, 16'hfff6, 16'h000d, 16'h000c, 16'h000f, 16'h0008, 16'h0000, 16'h0010, 16'hfff4, 16'hfffe, 16'hfff3, 16'hfff2, 16'h000b, 16'h0009, 16'hfff2, 16'h0001, 16'h000b, 16'h0010, 16'hfffb, 16'h0002, 16'hfffe, 16'h0003, 16'h000f, 16'h000d, 16'h0002, 16'hfff9, 16'hfff9, 16'h0009, 16'hfff7, 16'h000e, 16'h0002, 16'hfffc, 16'h0004, 16'hfff7, 16'hfff5, 16'hfffd, 16'h0001, 16'h0004, 16'h000b, 16'h0005, 16'h0002, 16'h0007, 16'hfff9, 16'hfff2, 16'h0006, 16'h000e, 16'h000b, 16'h0001, 16'h0004, 16'h000e, 16'h000b, 16'h0004, 16'h000c, 16'hffff, 16'h0000, 16'hfff4, 16'hfff1, 16'h0005, 16'hfff4, 16'hfff1, 16'h0002, 16'hfff6, 16'hfff5, 16'h000d, 16'h0008, 16'h0008, 16'h000e, 16'h0010 };
assign dw_3[3] = dw_3_3[d3_cntr];
