localparam D1_IN_SIZE = 1;
localparam D1_BW_W = 2;
localparam D1_SHIFT = 0;
localparam LOG2_D1_CYC = 9;
localparam D1_CYC = 512;
localparam D1_CH = 128;
reg [LOG2_D1_CYC-1:0] d1_cntr;
wire [D1_CH-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1;
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_0 = { 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3 };
assign dw_1[0] = dw_1_0[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_1 = { 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0 };
assign dw_1[1] = dw_1_1[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_2 = { 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1 };
assign dw_1[2] = dw_1_2[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_3 = { 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0 };
assign dw_1[3] = dw_1_3[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_4 = { 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3 };
assign dw_1[4] = dw_1_4[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_5 = { 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0 };
assign dw_1[5] = dw_1_5[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_6 = { 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3 };
assign dw_1[6] = dw_1_6[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_7 = { 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1 };
assign dw_1[7] = dw_1_7[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_8 = { 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1 };
assign dw_1[8] = dw_1_8[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_9 = { 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3 };
assign dw_1[9] = dw_1_9[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_10 = { 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3 };
assign dw_1[10] = dw_1_10[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_11 = { 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1 };
assign dw_1[11] = dw_1_11[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_12 = { 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3 };
assign dw_1[12] = dw_1_12[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_13 = { 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1 };
assign dw_1[13] = dw_1_13[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_14 = { 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3 };
assign dw_1[14] = dw_1_14[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_15 = { 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1 };
assign dw_1[15] = dw_1_15[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_16 = { 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0 };
assign dw_1[16] = dw_1_16[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_17 = { 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0 };
assign dw_1[17] = dw_1_17[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_18 = { 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0 };
assign dw_1[18] = dw_1_18[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_19 = { 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0 };
assign dw_1[19] = dw_1_19[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_20 = { 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0 };
assign dw_1[20] = dw_1_20[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_21 = { 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0 };
assign dw_1[21] = dw_1_21[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_22 = { 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1 };
assign dw_1[22] = dw_1_22[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_23 = { 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3 };
assign dw_1[23] = dw_1_23[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_24 = { 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3 };
assign dw_1[24] = dw_1_24[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_25 = { 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1 };
assign dw_1[25] = dw_1_25[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_26 = { 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3 };
assign dw_1[26] = dw_1_26[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_27 = { 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0 };
assign dw_1[27] = dw_1_27[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_28 = { 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1 };
assign dw_1[28] = dw_1_28[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_29 = { 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3 };
assign dw_1[29] = dw_1_29[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_30 = { 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0 };
assign dw_1[30] = dw_1_30[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_31 = { 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0 };
assign dw_1[31] = dw_1_31[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_32 = { 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0 };
assign dw_1[32] = dw_1_32[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_33 = { 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0 };
assign dw_1[33] = dw_1_33[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_34 = { 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0 };
assign dw_1[34] = dw_1_34[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_35 = { 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0 };
assign dw_1[35] = dw_1_35[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_36 = { 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1 };
assign dw_1[36] = dw_1_36[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_37 = { 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1 };
assign dw_1[37] = dw_1_37[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_38 = { 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1 };
assign dw_1[38] = dw_1_38[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_39 = { 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1 };
assign dw_1[39] = dw_1_39[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_40 = { 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1 };
assign dw_1[40] = dw_1_40[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_41 = { 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1 };
assign dw_1[41] = dw_1_41[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_42 = { 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0 };
assign dw_1[42] = dw_1_42[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_43 = { 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3 };
assign dw_1[43] = dw_1_43[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_44 = { 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0 };
assign dw_1[44] = dw_1_44[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_45 = { 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3 };
assign dw_1[45] = dw_1_45[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_46 = { 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0 };
assign dw_1[46] = dw_1_46[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_47 = { 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3 };
assign dw_1[47] = dw_1_47[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_48 = { 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0 };
assign dw_1[48] = dw_1_48[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_49 = { 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0 };
assign dw_1[49] = dw_1_49[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_50 = { 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1 };
assign dw_1[50] = dw_1_50[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_51 = { 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0 };
assign dw_1[51] = dw_1_51[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_52 = { 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3 };
assign dw_1[52] = dw_1_52[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_53 = { 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1 };
assign dw_1[53] = dw_1_53[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_54 = { 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0 };
assign dw_1[54] = dw_1_54[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_55 = { 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0 };
assign dw_1[55] = dw_1_55[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_56 = { 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1 };
assign dw_1[56] = dw_1_56[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_57 = { 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3 };
assign dw_1[57] = dw_1_57[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_58 = { 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1 };
assign dw_1[58] = dw_1_58[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_59 = { 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3 };
assign dw_1[59] = dw_1_59[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_60 = { 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0 };
assign dw_1[60] = dw_1_60[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_61 = { 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0 };
assign dw_1[61] = dw_1_61[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_62 = { 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0 };
assign dw_1[62] = dw_1_62[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_63 = { 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3 };
assign dw_1[63] = dw_1_63[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_64 = { 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3 };
assign dw_1[64] = dw_1_64[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_65 = { 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3 };
assign dw_1[65] = dw_1_65[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_66 = { 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3 };
assign dw_1[66] = dw_1_66[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_67 = { 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1 };
assign dw_1[67] = dw_1_67[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_68 = { 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3 };
assign dw_1[68] = dw_1_68[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_69 = { 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0 };
assign dw_1[69] = dw_1_69[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_70 = { 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1 };
assign dw_1[70] = dw_1_70[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_71 = { 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1 };
assign dw_1[71] = dw_1_71[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_72 = { 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0 };
assign dw_1[72] = dw_1_72[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_73 = { 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3 };
assign dw_1[73] = dw_1_73[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_74 = { 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3 };
assign dw_1[74] = dw_1_74[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_75 = { 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3 };
assign dw_1[75] = dw_1_75[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_76 = { 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1 };
assign dw_1[76] = dw_1_76[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_77 = { 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0 };
assign dw_1[77] = dw_1_77[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_78 = { 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0 };
assign dw_1[78] = dw_1_78[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_79 = { 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0 };
assign dw_1[79] = dw_1_79[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_80 = { 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1 };
assign dw_1[80] = dw_1_80[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_81 = { 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3 };
assign dw_1[81] = dw_1_81[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_82 = { 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0 };
assign dw_1[82] = dw_1_82[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_83 = { 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3 };
assign dw_1[83] = dw_1_83[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_84 = { 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3 };
assign dw_1[84] = dw_1_84[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_85 = { 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3 };
assign dw_1[85] = dw_1_85[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_86 = { 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0 };
assign dw_1[86] = dw_1_86[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_87 = { 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0 };
assign dw_1[87] = dw_1_87[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_88 = { 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3 };
assign dw_1[88] = dw_1_88[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_89 = { 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0 };
assign dw_1[89] = dw_1_89[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_90 = { 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0 };
assign dw_1[90] = dw_1_90[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_91 = { 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0 };
assign dw_1[91] = dw_1_91[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_92 = { 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0 };
assign dw_1[92] = dw_1_92[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_93 = { 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3 };
assign dw_1[93] = dw_1_93[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_94 = { 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1 };
assign dw_1[94] = dw_1_94[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_95 = { 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1 };
assign dw_1[95] = dw_1_95[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_96 = { 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1 };
assign dw_1[96] = dw_1_96[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_97 = { 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3 };
assign dw_1[97] = dw_1_97[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_98 = { 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0 };
assign dw_1[98] = dw_1_98[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_99 = { 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1 };
assign dw_1[99] = dw_1_99[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_100 = { 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0 };
assign dw_1[100] = dw_1_100[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_101 = { 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0 };
assign dw_1[101] = dw_1_101[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_102 = { 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0 };
assign dw_1[102] = dw_1_102[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_103 = { 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1 };
assign dw_1[103] = dw_1_103[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_104 = { 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3 };
assign dw_1[104] = dw_1_104[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_105 = { 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1 };
assign dw_1[105] = dw_1_105[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_106 = { 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1 };
assign dw_1[106] = dw_1_106[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_107 = { 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3 };
assign dw_1[107] = dw_1_107[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_108 = { 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3 };
assign dw_1[108] = dw_1_108[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_109 = { 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0 };
assign dw_1[109] = dw_1_109[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_110 = { 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1 };
assign dw_1[110] = dw_1_110[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_111 = { 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3 };
assign dw_1[111] = dw_1_111[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_112 = { 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3 };
assign dw_1[112] = dw_1_112[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_113 = { 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3 };
assign dw_1[113] = dw_1_113[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_114 = { 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0 };
assign dw_1[114] = dw_1_114[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_115 = { 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3 };
assign dw_1[115] = dw_1_115[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_116 = { 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3 };
assign dw_1[116] = dw_1_116[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_117 = { 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0 };
assign dw_1[117] = dw_1_117[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_118 = { 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3 };
assign dw_1[118] = dw_1_118[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_119 = { 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3 };
assign dw_1[119] = dw_1_119[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_120 = { 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1 };
assign dw_1[120] = dw_1_120[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_121 = { 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0 };
assign dw_1[121] = dw_1_121[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_122 = { 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0 };
assign dw_1[122] = dw_1_122[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_123 = { 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0 };
assign dw_1[123] = dw_1_123[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_124 = { 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3 };
assign dw_1[124] = dw_1_124[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_125 = { 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1 };
assign dw_1[125] = dw_1_125[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_126 = { 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0 };
assign dw_1[126] = dw_1_126[d1_cntr];
reg [D1_CYC-1:0][D1_IN_SIZE*D1_BW_W-1:0] dw_1_127 = { 2'h1, 2'h0, 2'h1, 2'h0, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h1, 2'h1, 2'h1, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h1, 2'h3, 2'h1, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h1, 2'h1, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h0, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h1, 2'h0, 2'h1, 2'h3, 2'h0, 2'h0, 2'h3, 2'h1, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h1, 2'h0, 2'h1, 2'h1, 2'h0, 2'h1, 2'h3, 2'h3, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h0, 2'h3, 2'h0, 2'h3, 2'h0, 2'h0, 2'h1, 2'h1, 2'h3, 2'h3, 2'h3, 2'h0, 2'h0, 2'h3, 2'h3, 2'h3, 2'h0, 2'h3, 2'h3, 2'h1, 2'h1, 2'h0, 2'h0, 2'h0, 2'h0, 2'h0, 2'h1, 2'h3, 2'h1, 2'h0, 2'h1, 2'h0, 2'h0, 2'h1, 2'h3, 2'h0, 2'h3, 2'h3, 2'h0, 2'h3 };
assign dw_1[127] = dw_1_127[d1_cntr];
